magic
tech sky130A
magscale 1 2
timestamp 1748334013
<< metal1 >>
rect 0 44952 200 45152
rect 28872 44952 29072 45152
rect 21549 41418 21601 41424
rect 21549 41360 21601 41366
rect 21849 41418 21901 41424
rect 21849 41360 21901 41366
rect 22149 41418 22201 41424
rect 22149 41360 22201 41366
rect 22449 41418 22501 41424
rect 22449 41360 22501 41366
rect 22749 41418 22801 41424
rect 22749 41360 22801 41366
rect 23049 41418 23101 41424
rect 23049 41360 23101 41366
rect 23349 41418 23401 41424
rect 23349 41360 23401 41366
rect 23649 41418 23701 41424
rect 23649 41360 23701 41366
rect 3933 40630 3985 40636
rect 3933 40572 3985 40578
rect 4233 40630 4285 40636
rect 4233 40572 4285 40578
rect 4533 40630 4585 40636
rect 4533 40572 4585 40578
rect 4833 40630 4885 40636
rect 4833 40572 4885 40578
rect 5133 40630 5185 40636
rect 5133 40572 5185 40578
rect 5433 40630 5485 40636
rect 5433 40572 5485 40578
rect 5733 40630 5785 40636
rect 5733 40572 5785 40578
rect 6033 40630 6085 40636
rect 6033 40572 6085 40578
rect 8349 40630 8401 40636
rect 8349 40572 8401 40578
rect 8649 40630 8701 40636
rect 8649 40572 8701 40578
rect 8949 40630 9001 40636
rect 8949 40572 9001 40578
rect 9249 40630 9301 40636
rect 9249 40572 9301 40578
rect 9549 40630 9601 40636
rect 9549 40572 9601 40578
rect 9849 40630 9901 40636
rect 9849 40572 9901 40578
rect 10149 40630 10201 40636
rect 10149 40572 10201 40578
rect 10449 40630 10501 40636
rect 10449 40572 10501 40578
rect 12765 40630 12817 40636
rect 12765 40572 12817 40578
rect 13065 40630 13117 40636
rect 13065 40572 13117 40578
rect 13365 40630 13417 40636
rect 13365 40572 13417 40578
rect 13665 40630 13717 40636
rect 13665 40572 13717 40578
rect 13965 40630 14017 40636
rect 13965 40572 14017 40578
rect 14265 40630 14317 40636
rect 14265 40572 14317 40578
rect 14565 40630 14617 40636
rect 14565 40572 14617 40578
rect 14865 40630 14917 40636
rect 14865 40572 14917 40578
rect 21640 37862 21692 37868
rect 21640 37804 21692 37810
rect 21940 37862 21992 37868
rect 21940 37804 21992 37810
rect 22240 37862 22292 37868
rect 22240 37804 22292 37810
rect 22540 37862 22592 37868
rect 22540 37804 22592 37810
rect 22840 37862 22892 37868
rect 22840 37804 22892 37810
rect 23140 37862 23192 37868
rect 23140 37804 23192 37810
rect 23440 37862 23492 37868
rect 23440 37804 23492 37810
rect 23740 37862 23792 37868
rect 23740 37804 23792 37810
rect 0 0 200 200
rect 28872 0 29072 200
<< via1 >>
rect 21549 41366 21601 41418
rect 21849 41366 21901 41418
rect 22149 41366 22201 41418
rect 22449 41366 22501 41418
rect 22749 41366 22801 41418
rect 23049 41366 23101 41418
rect 23349 41366 23401 41418
rect 23649 41366 23701 41418
rect 3933 40578 3985 40630
rect 4233 40578 4285 40630
rect 4533 40578 4585 40630
rect 4833 40578 4885 40630
rect 5133 40578 5185 40630
rect 5433 40578 5485 40630
rect 5733 40578 5785 40630
rect 6033 40578 6085 40630
rect 8349 40578 8401 40630
rect 8649 40578 8701 40630
rect 8949 40578 9001 40630
rect 9249 40578 9301 40630
rect 9549 40578 9601 40630
rect 9849 40578 9901 40630
rect 10149 40578 10201 40630
rect 10449 40578 10501 40630
rect 12765 40578 12817 40630
rect 13065 40578 13117 40630
rect 13365 40578 13417 40630
rect 13665 40578 13717 40630
rect 13965 40578 14017 40630
rect 14265 40578 14317 40630
rect 14565 40578 14617 40630
rect 14865 40578 14917 40630
rect 21640 37810 21692 37862
rect 21940 37810 21992 37862
rect 22240 37810 22292 37862
rect 22540 37810 22592 37862
rect 22840 37810 22892 37862
rect 23140 37810 23192 37862
rect 23440 37810 23492 37862
rect 23740 37810 23792 37862
<< metal2 >>
rect 3520 39679 3620 41576
rect 3670 40384 3770 41576
rect 3931 40632 3987 40641
rect 4231 40632 4287 40641
rect 4531 40632 4587 40641
rect 4831 40632 4887 40641
rect 5131 40632 5187 40641
rect 5431 40632 5487 40641
rect 5731 40632 5787 40641
rect 6031 40632 6087 40641
rect 3927 40578 3931 40630
rect 3987 40578 3991 40630
rect 4227 40578 4231 40630
rect 4287 40578 4291 40630
rect 4527 40578 4531 40630
rect 4587 40578 4591 40630
rect 4827 40578 4831 40630
rect 4887 40578 4891 40630
rect 5127 40578 5131 40630
rect 5187 40578 5191 40630
rect 5427 40578 5431 40630
rect 5487 40578 5491 40630
rect 5727 40578 5731 40630
rect 5787 40578 5791 40630
rect 6027 40578 6031 40630
rect 6087 40578 6091 40630
rect 3931 40567 3987 40576
rect 4231 40567 4287 40576
rect 4531 40567 4587 40576
rect 4831 40567 4887 40576
rect 5131 40567 5187 40576
rect 5431 40567 5487 40576
rect 5731 40567 5787 40576
rect 6031 40567 6087 40576
rect 6166 40384 6266 41576
rect 3670 40284 3870 40384
rect 3770 40079 3870 40284
rect 6066 40284 6266 40384
rect 6066 40079 6166 40284
rect 3716 39889 3725 40079
rect 3915 39889 3924 40079
rect 6012 39889 6021 40079
rect 6211 39889 6220 40079
rect 6316 39679 6416 41576
rect 7936 39679 8036 41576
rect 8086 40384 8186 41576
rect 8347 40632 8403 40641
rect 8647 40632 8703 40641
rect 8947 40632 9003 40641
rect 9247 40632 9303 40641
rect 9547 40632 9603 40641
rect 9847 40632 9903 40641
rect 10147 40632 10203 40641
rect 10447 40632 10503 40641
rect 8343 40578 8347 40630
rect 8403 40578 8407 40630
rect 8643 40578 8647 40630
rect 8703 40578 8707 40630
rect 8943 40578 8947 40630
rect 9003 40578 9007 40630
rect 9243 40578 9247 40630
rect 9303 40578 9307 40630
rect 9543 40578 9547 40630
rect 9603 40578 9607 40630
rect 9843 40578 9847 40630
rect 9903 40578 9907 40630
rect 10143 40578 10147 40630
rect 10203 40578 10207 40630
rect 10443 40578 10447 40630
rect 10503 40578 10507 40630
rect 8347 40567 8403 40576
rect 8647 40567 8703 40576
rect 8947 40567 9003 40576
rect 9247 40567 9303 40576
rect 9547 40567 9603 40576
rect 9847 40567 9903 40576
rect 10147 40567 10203 40576
rect 10447 40567 10503 40576
rect 10582 40384 10682 41576
rect 8086 40284 8286 40384
rect 8186 40079 8286 40284
rect 10482 40284 10682 40384
rect 10482 40079 10582 40284
rect 8132 39889 8141 40079
rect 8331 39889 8340 40079
rect 10428 39889 10437 40079
rect 10627 39889 10636 40079
rect 10732 39679 10832 41576
rect 12352 39679 12452 41576
rect 12502 40384 12602 41576
rect 12763 40632 12819 40641
rect 13063 40632 13119 40641
rect 13363 40632 13419 40641
rect 13663 40632 13719 40641
rect 13963 40632 14019 40641
rect 14263 40632 14319 40641
rect 14563 40632 14619 40641
rect 14863 40632 14919 40641
rect 12759 40578 12763 40630
rect 12819 40578 12823 40630
rect 13059 40578 13063 40630
rect 13119 40578 13123 40630
rect 13359 40578 13363 40630
rect 13419 40578 13423 40630
rect 13659 40578 13663 40630
rect 13719 40578 13723 40630
rect 13959 40578 13963 40630
rect 14019 40578 14023 40630
rect 14259 40578 14263 40630
rect 14319 40578 14323 40630
rect 14559 40578 14563 40630
rect 14619 40578 14623 40630
rect 14859 40578 14863 40630
rect 14919 40578 14923 40630
rect 12763 40567 12819 40576
rect 13063 40567 13119 40576
rect 13363 40567 13419 40576
rect 13663 40567 13719 40576
rect 13963 40567 14019 40576
rect 14263 40567 14319 40576
rect 14563 40567 14619 40576
rect 14863 40567 14919 40576
rect 14998 40384 15098 41576
rect 12502 40284 12702 40384
rect 12602 40079 12702 40284
rect 14898 40284 15098 40384
rect 14898 40079 14998 40284
rect 12548 39889 12557 40079
rect 12747 39889 12756 40079
rect 14844 39889 14853 40079
rect 15043 39889 15052 40079
rect 15148 39679 15248 41576
rect 21547 41420 21603 41429
rect 21847 41420 21903 41429
rect 22147 41420 22203 41429
rect 22447 41420 22503 41429
rect 22747 41420 22803 41429
rect 23047 41420 23103 41429
rect 23347 41420 23403 41429
rect 23647 41420 23703 41429
rect 21543 41366 21547 41418
rect 21603 41366 21607 41418
rect 21843 41366 21847 41418
rect 21903 41366 21907 41418
rect 22143 41366 22147 41418
rect 22203 41366 22207 41418
rect 22443 41366 22447 41418
rect 22503 41366 22507 41418
rect 22743 41366 22747 41418
rect 22803 41366 22807 41418
rect 23043 41366 23047 41418
rect 23103 41366 23107 41418
rect 23343 41366 23347 41418
rect 23403 41366 23407 41418
rect 23643 41366 23647 41418
rect 23703 41366 23707 41418
rect 21547 41355 21603 41364
rect 21847 41355 21903 41364
rect 22147 41355 22203 41364
rect 22447 41355 22503 41364
rect 22747 41355 22803 41364
rect 23047 41355 23103 41364
rect 23347 41355 23403 41364
rect 23647 41355 23703 41364
rect 21274 40684 21284 40884
rect 21474 40684 21483 40884
rect 23780 40684 23789 40884
rect 23979 40684 23989 40884
rect 21024 40284 21034 40484
rect 21224 40284 21233 40484
rect 24030 40284 24039 40484
rect 24229 40284 24239 40484
rect 21274 39884 21284 40084
rect 21474 39884 21483 40084
rect 3466 39489 3475 39679
rect 3665 39489 3674 39679
rect 6262 39489 6271 39679
rect 6461 39489 6470 39679
rect 7882 39489 7891 39679
rect 8081 39489 8090 39679
rect 10678 39489 10687 39679
rect 10877 39489 10886 39679
rect 12298 39489 12307 39679
rect 12497 39489 12506 39679
rect 15094 39489 15103 39679
rect 15293 39489 15302 39679
rect 23780 38284 23789 38484
rect 23979 38284 23989 38484
rect 21638 37864 21694 37873
rect 21938 37864 21994 37873
rect 22238 37864 22294 37873
rect 22538 37864 22594 37873
rect 22838 37864 22894 37873
rect 23138 37864 23194 37873
rect 23438 37864 23494 37873
rect 23738 37864 23794 37873
rect 21634 37810 21638 37862
rect 21694 37810 21698 37862
rect 21934 37810 21938 37862
rect 21994 37810 21998 37862
rect 22234 37810 22238 37862
rect 22294 37810 22298 37862
rect 22534 37810 22538 37862
rect 22594 37810 22598 37862
rect 22834 37810 22838 37862
rect 22894 37810 22898 37862
rect 23134 37810 23138 37862
rect 23194 37810 23198 37862
rect 23434 37810 23438 37862
rect 23494 37810 23498 37862
rect 23734 37810 23738 37862
rect 23794 37810 23798 37862
rect 21638 37799 21694 37808
rect 21938 37799 21994 37808
rect 22238 37799 22294 37808
rect 22538 37799 22594 37808
rect 22838 37799 22894 37808
rect 23138 37799 23194 37808
rect 23438 37799 23494 37808
rect 23738 37799 23794 37808
rect 21507 26103 21677 26107
rect 23018 26103 23188 26107
rect 21502 26098 23193 26103
rect 21502 25928 21507 26098
rect 21677 25928 23018 26098
rect 23188 25928 23193 26098
rect 21502 25923 23193 25928
rect 21507 25919 21677 25923
rect 23018 25919 23188 25923
<< via2 >>
rect 3931 40630 3987 40632
rect 4231 40630 4287 40632
rect 4531 40630 4587 40632
rect 4831 40630 4887 40632
rect 5131 40630 5187 40632
rect 5431 40630 5487 40632
rect 5731 40630 5787 40632
rect 6031 40630 6087 40632
rect 3931 40578 3933 40630
rect 3933 40578 3985 40630
rect 3985 40578 3987 40630
rect 4231 40578 4233 40630
rect 4233 40578 4285 40630
rect 4285 40578 4287 40630
rect 4531 40578 4533 40630
rect 4533 40578 4585 40630
rect 4585 40578 4587 40630
rect 4831 40578 4833 40630
rect 4833 40578 4885 40630
rect 4885 40578 4887 40630
rect 5131 40578 5133 40630
rect 5133 40578 5185 40630
rect 5185 40578 5187 40630
rect 5431 40578 5433 40630
rect 5433 40578 5485 40630
rect 5485 40578 5487 40630
rect 5731 40578 5733 40630
rect 5733 40578 5785 40630
rect 5785 40578 5787 40630
rect 6031 40578 6033 40630
rect 6033 40578 6085 40630
rect 6085 40578 6087 40630
rect 3931 40576 3987 40578
rect 4231 40576 4287 40578
rect 4531 40576 4587 40578
rect 4831 40576 4887 40578
rect 5131 40576 5187 40578
rect 5431 40576 5487 40578
rect 5731 40576 5787 40578
rect 6031 40576 6087 40578
rect 3725 39889 3915 40079
rect 6021 39889 6211 40079
rect 8347 40630 8403 40632
rect 8647 40630 8703 40632
rect 8947 40630 9003 40632
rect 9247 40630 9303 40632
rect 9547 40630 9603 40632
rect 9847 40630 9903 40632
rect 10147 40630 10203 40632
rect 10447 40630 10503 40632
rect 8347 40578 8349 40630
rect 8349 40578 8401 40630
rect 8401 40578 8403 40630
rect 8647 40578 8649 40630
rect 8649 40578 8701 40630
rect 8701 40578 8703 40630
rect 8947 40578 8949 40630
rect 8949 40578 9001 40630
rect 9001 40578 9003 40630
rect 9247 40578 9249 40630
rect 9249 40578 9301 40630
rect 9301 40578 9303 40630
rect 9547 40578 9549 40630
rect 9549 40578 9601 40630
rect 9601 40578 9603 40630
rect 9847 40578 9849 40630
rect 9849 40578 9901 40630
rect 9901 40578 9903 40630
rect 10147 40578 10149 40630
rect 10149 40578 10201 40630
rect 10201 40578 10203 40630
rect 10447 40578 10449 40630
rect 10449 40578 10501 40630
rect 10501 40578 10503 40630
rect 8347 40576 8403 40578
rect 8647 40576 8703 40578
rect 8947 40576 9003 40578
rect 9247 40576 9303 40578
rect 9547 40576 9603 40578
rect 9847 40576 9903 40578
rect 10147 40576 10203 40578
rect 10447 40576 10503 40578
rect 8141 39889 8331 40079
rect 10437 39889 10627 40079
rect 12763 40630 12819 40632
rect 13063 40630 13119 40632
rect 13363 40630 13419 40632
rect 13663 40630 13719 40632
rect 13963 40630 14019 40632
rect 14263 40630 14319 40632
rect 14563 40630 14619 40632
rect 14863 40630 14919 40632
rect 12763 40578 12765 40630
rect 12765 40578 12817 40630
rect 12817 40578 12819 40630
rect 13063 40578 13065 40630
rect 13065 40578 13117 40630
rect 13117 40578 13119 40630
rect 13363 40578 13365 40630
rect 13365 40578 13417 40630
rect 13417 40578 13419 40630
rect 13663 40578 13665 40630
rect 13665 40578 13717 40630
rect 13717 40578 13719 40630
rect 13963 40578 13965 40630
rect 13965 40578 14017 40630
rect 14017 40578 14019 40630
rect 14263 40578 14265 40630
rect 14265 40578 14317 40630
rect 14317 40578 14319 40630
rect 14563 40578 14565 40630
rect 14565 40578 14617 40630
rect 14617 40578 14619 40630
rect 14863 40578 14865 40630
rect 14865 40578 14917 40630
rect 14917 40578 14919 40630
rect 12763 40576 12819 40578
rect 13063 40576 13119 40578
rect 13363 40576 13419 40578
rect 13663 40576 13719 40578
rect 13963 40576 14019 40578
rect 14263 40576 14319 40578
rect 14563 40576 14619 40578
rect 14863 40576 14919 40578
rect 12557 39889 12747 40079
rect 14853 39889 15043 40079
rect 21547 41418 21603 41420
rect 21847 41418 21903 41420
rect 22147 41418 22203 41420
rect 22447 41418 22503 41420
rect 22747 41418 22803 41420
rect 23047 41418 23103 41420
rect 23347 41418 23403 41420
rect 23647 41418 23703 41420
rect 21547 41366 21549 41418
rect 21549 41366 21601 41418
rect 21601 41366 21603 41418
rect 21847 41366 21849 41418
rect 21849 41366 21901 41418
rect 21901 41366 21903 41418
rect 22147 41366 22149 41418
rect 22149 41366 22201 41418
rect 22201 41366 22203 41418
rect 22447 41366 22449 41418
rect 22449 41366 22501 41418
rect 22501 41366 22503 41418
rect 22747 41366 22749 41418
rect 22749 41366 22801 41418
rect 22801 41366 22803 41418
rect 23047 41366 23049 41418
rect 23049 41366 23101 41418
rect 23101 41366 23103 41418
rect 23347 41366 23349 41418
rect 23349 41366 23401 41418
rect 23401 41366 23403 41418
rect 23647 41366 23649 41418
rect 23649 41366 23701 41418
rect 23701 41366 23703 41418
rect 21547 41364 21603 41366
rect 21847 41364 21903 41366
rect 22147 41364 22203 41366
rect 22447 41364 22503 41366
rect 22747 41364 22803 41366
rect 23047 41364 23103 41366
rect 23347 41364 23403 41366
rect 23647 41364 23703 41366
rect 21284 40684 21474 40884
rect 23789 40684 23979 40884
rect 21034 40284 21224 40484
rect 24039 40284 24229 40484
rect 21284 39884 21474 40084
rect 3475 39489 3665 39679
rect 6271 39489 6461 39679
rect 7891 39489 8081 39679
rect 10687 39489 10877 39679
rect 12307 39489 12497 39679
rect 15103 39489 15293 39679
rect 23789 38284 23979 38484
rect 21638 37862 21694 37864
rect 21938 37862 21994 37864
rect 22238 37862 22294 37864
rect 22538 37862 22594 37864
rect 22838 37862 22894 37864
rect 23138 37862 23194 37864
rect 23438 37862 23494 37864
rect 23738 37862 23794 37864
rect 21638 37810 21640 37862
rect 21640 37810 21692 37862
rect 21692 37810 21694 37862
rect 21938 37810 21940 37862
rect 21940 37810 21992 37862
rect 21992 37810 21994 37862
rect 22238 37810 22240 37862
rect 22240 37810 22292 37862
rect 22292 37810 22294 37862
rect 22538 37810 22540 37862
rect 22540 37810 22592 37862
rect 22592 37810 22594 37862
rect 22838 37810 22840 37862
rect 22840 37810 22892 37862
rect 22892 37810 22894 37862
rect 23138 37810 23140 37862
rect 23140 37810 23192 37862
rect 23192 37810 23194 37862
rect 23438 37810 23440 37862
rect 23440 37810 23492 37862
rect 23492 37810 23494 37862
rect 23738 37810 23740 37862
rect 23740 37810 23792 37862
rect 23792 37810 23794 37862
rect 21638 37808 21694 37810
rect 21938 37808 21994 37810
rect 22238 37808 22294 37810
rect 22538 37808 22594 37810
rect 22838 37808 22894 37810
rect 23138 37808 23194 37810
rect 23438 37808 23494 37810
rect 23738 37808 23794 37810
rect 21507 25928 21677 26098
rect 23018 25928 23188 26098
<< metal3 >>
rect 2998 44950 3004 45014
rect 3068 44950 3074 45014
rect 3550 44950 3556 45014
rect 3620 44950 3626 45014
rect 4102 44950 4108 45014
rect 4172 44950 4178 45014
rect 4654 44950 4660 45014
rect 4724 44950 4730 45014
rect 5206 44950 5212 45014
rect 5276 44950 5282 45014
rect 5758 44950 5764 45014
rect 5828 44950 5834 45014
rect 6310 44950 6316 45014
rect 6380 44950 6386 45014
rect 6862 44950 6868 45014
rect 6932 44950 6938 45014
rect 7414 44950 7420 45014
rect 7484 44950 7490 45014
rect 7966 44950 7972 45014
rect 8036 44950 8042 45014
rect 8518 44950 8524 45014
rect 8588 44950 8594 45014
rect 9070 44950 9076 45014
rect 9140 44950 9146 45014
rect 9622 44950 9628 45014
rect 9692 44950 9698 45014
rect 10174 44950 10180 45014
rect 10244 44950 10250 45014
rect 10726 44950 10732 45014
rect 10796 44950 10802 45014
rect 11278 44950 11284 45014
rect 11348 44950 11354 45014
rect 11830 44950 11836 45014
rect 11900 44950 11906 45014
rect 12382 44950 12388 45014
rect 12452 44950 12458 45014
rect 12934 44950 12940 45014
rect 13004 44950 13010 45014
rect 13486 44950 13492 45014
rect 13556 44950 13562 45014
rect 14038 44950 14044 45014
rect 14108 44950 14114 45014
rect 14590 44950 14596 45014
rect 14660 44950 14666 45014
rect 15142 44950 15148 45014
rect 15212 44950 15218 45014
rect 15694 44950 15700 45014
rect 15764 44950 15770 45014
rect 20662 44950 20668 45014
rect 20732 44950 20738 45014
rect 21214 44950 21220 45014
rect 21284 44950 21290 45014
rect 21766 44950 21772 45014
rect 21836 44950 21842 45014
rect 22318 44950 22324 45014
rect 22388 44950 22394 45014
rect 22870 44950 22876 45014
rect 22940 44950 22946 45014
rect 23422 44950 23428 45014
rect 23492 44950 23498 45014
rect 23974 44952 23980 45016
rect 24044 44952 24050 45016
rect 3006 41776 3066 44950
rect 3558 41976 3618 44950
rect 4110 42176 4170 44950
rect 4662 42376 4722 44950
rect 5214 42376 5274 44950
rect 4662 42316 4889 42376
rect 4110 42116 4589 42176
rect 3558 41916 4289 41976
rect 3006 41716 3989 41776
rect 3929 40637 3989 41716
rect 4229 40637 4289 41916
rect 4529 40637 4589 42116
rect 4829 40637 4889 42316
rect 5129 42316 5274 42376
rect 5129 40637 5189 42316
rect 5766 42176 5826 44950
rect 5429 42116 5826 42176
rect 5429 40637 5489 42116
rect 6318 41976 6378 44950
rect 5729 41916 6378 41976
rect 5729 40637 5789 41916
rect 6870 41776 6930 44950
rect 6029 41716 6930 41776
rect 7422 41776 7482 44950
rect 7974 41976 8034 44950
rect 8526 42176 8586 44950
rect 9078 42376 9138 44950
rect 9630 42376 9690 44950
rect 9078 42316 9305 42376
rect 8526 42116 9005 42176
rect 7974 41916 8705 41976
rect 7422 41716 8405 41776
rect 6029 40637 6089 41716
rect 8345 40637 8405 41716
rect 8645 40637 8705 41916
rect 8945 40637 9005 42116
rect 9245 40637 9305 42316
rect 9545 42316 9690 42376
rect 9545 40637 9605 42316
rect 10182 42176 10242 44950
rect 9845 42116 10242 42176
rect 9845 40637 9905 42116
rect 10734 41976 10794 44950
rect 10145 41916 10794 41976
rect 10145 40637 10205 41916
rect 11286 41776 11346 44950
rect 10445 41716 11346 41776
rect 11838 41776 11898 44950
rect 12390 41976 12450 44950
rect 12942 42176 13002 44950
rect 13494 42376 13554 44950
rect 14046 42376 14106 44950
rect 13494 42316 13721 42376
rect 12942 42116 13421 42176
rect 12390 41916 13121 41976
rect 11838 41716 12821 41776
rect 10445 40637 10505 41716
rect 12761 40637 12821 41716
rect 13061 40637 13121 41916
rect 13361 40637 13421 42116
rect 13661 40637 13721 42316
rect 13961 42316 14106 42376
rect 13961 40637 14021 42316
rect 14598 42176 14658 44950
rect 14261 42116 14658 42176
rect 14261 40637 14321 42116
rect 15150 41976 15210 44950
rect 14561 41916 15210 41976
rect 14561 40637 14621 41916
rect 15702 41776 15762 44950
rect 14861 41716 15762 41776
rect 20670 41775 20730 44950
rect 21222 41975 21282 44950
rect 21774 42175 21834 44950
rect 22326 42372 22386 44950
rect 22878 42375 22938 44950
rect 22326 42312 22505 42372
rect 21774 42115 22205 42175
rect 21222 41915 21905 41975
rect 14861 40637 14921 41716
rect 20670 41715 21605 41775
rect 21545 41425 21605 41715
rect 21845 41425 21905 41915
rect 22145 41425 22205 42115
rect 22445 41425 22505 42312
rect 22745 42315 22938 42375
rect 22745 41425 22805 42315
rect 23430 42175 23490 44950
rect 23045 42115 23490 42175
rect 23045 41425 23105 42115
rect 23982 41975 24042 44952
rect 24526 44950 24532 45014
rect 24596 44950 24602 45014
rect 23345 41915 24042 41975
rect 23345 41425 23405 41915
rect 24534 41775 24594 44950
rect 23645 41715 24594 41775
rect 23645 41425 23705 41715
rect 21542 41420 21608 41425
rect 21542 41364 21547 41420
rect 21603 41364 21608 41420
rect 21542 41359 21608 41364
rect 21842 41420 21908 41425
rect 21842 41364 21847 41420
rect 21903 41364 21908 41420
rect 21842 41359 21908 41364
rect 22142 41420 22208 41425
rect 22142 41364 22147 41420
rect 22203 41364 22208 41420
rect 22142 41359 22208 41364
rect 22442 41420 22508 41425
rect 22442 41364 22447 41420
rect 22503 41364 22508 41420
rect 22442 41359 22508 41364
rect 22742 41420 22808 41425
rect 22742 41364 22747 41420
rect 22803 41364 22808 41420
rect 22742 41359 22808 41364
rect 23042 41420 23108 41425
rect 23042 41364 23047 41420
rect 23103 41364 23108 41420
rect 23042 41359 23108 41364
rect 23342 41420 23408 41425
rect 23342 41364 23347 41420
rect 23403 41364 23408 41420
rect 23342 41359 23408 41364
rect 23642 41420 23708 41425
rect 23642 41364 23647 41420
rect 23703 41364 23708 41420
rect 23642 41359 23708 41364
rect 19700 40884 19900 40890
rect 21279 40884 21479 40889
rect 23784 40884 23984 40889
rect 19900 40686 21284 40884
rect 19700 40684 21284 40686
rect 21474 40684 23789 40884
rect 23979 40684 24139 40884
rect 19700 40680 19900 40684
rect 21279 40679 21479 40684
rect 23784 40679 23984 40684
rect 3926 40632 3992 40637
rect 3926 40576 3931 40632
rect 3987 40576 3992 40632
rect 3926 40571 3992 40576
rect 4226 40632 4292 40637
rect 4226 40576 4231 40632
rect 4287 40576 4292 40632
rect 4226 40571 4292 40576
rect 4526 40632 4592 40637
rect 4526 40576 4531 40632
rect 4587 40576 4592 40632
rect 4526 40571 4592 40576
rect 4826 40632 4892 40637
rect 4826 40576 4831 40632
rect 4887 40576 4892 40632
rect 4826 40571 4892 40576
rect 5126 40632 5192 40637
rect 5126 40576 5131 40632
rect 5187 40576 5192 40632
rect 5126 40571 5192 40576
rect 5426 40632 5492 40637
rect 5426 40576 5431 40632
rect 5487 40576 5492 40632
rect 5426 40571 5492 40576
rect 5726 40632 5792 40637
rect 5726 40576 5731 40632
rect 5787 40576 5792 40632
rect 5726 40571 5792 40576
rect 6026 40632 6092 40637
rect 6026 40576 6031 40632
rect 6087 40576 6092 40632
rect 6026 40571 6092 40576
rect 8342 40632 8408 40637
rect 8342 40576 8347 40632
rect 8403 40576 8408 40632
rect 8342 40571 8408 40576
rect 8642 40632 8708 40637
rect 8642 40576 8647 40632
rect 8703 40576 8708 40632
rect 8642 40571 8708 40576
rect 8942 40632 9008 40637
rect 8942 40576 8947 40632
rect 9003 40576 9008 40632
rect 8942 40571 9008 40576
rect 9242 40632 9308 40637
rect 9242 40576 9247 40632
rect 9303 40576 9308 40632
rect 9242 40571 9308 40576
rect 9542 40632 9608 40637
rect 9542 40576 9547 40632
rect 9603 40576 9608 40632
rect 9542 40571 9608 40576
rect 9842 40632 9908 40637
rect 9842 40576 9847 40632
rect 9903 40576 9908 40632
rect 9842 40571 9908 40576
rect 10142 40632 10208 40637
rect 10142 40576 10147 40632
rect 10203 40576 10208 40632
rect 10142 40571 10208 40576
rect 10442 40632 10508 40637
rect 10442 40576 10447 40632
rect 10503 40576 10508 40632
rect 10442 40571 10508 40576
rect 12758 40632 12824 40637
rect 12758 40576 12763 40632
rect 12819 40576 12824 40632
rect 12758 40571 12824 40576
rect 13058 40632 13124 40637
rect 13058 40576 13063 40632
rect 13119 40576 13124 40632
rect 13058 40571 13124 40576
rect 13358 40632 13424 40637
rect 13358 40576 13363 40632
rect 13419 40576 13424 40632
rect 13358 40571 13424 40576
rect 13658 40632 13724 40637
rect 13658 40576 13663 40632
rect 13719 40576 13724 40632
rect 13658 40571 13724 40576
rect 13958 40632 14024 40637
rect 13958 40576 13963 40632
rect 14019 40576 14024 40632
rect 13958 40571 14024 40576
rect 14258 40632 14324 40637
rect 14258 40576 14263 40632
rect 14319 40576 14324 40632
rect 14258 40571 14324 40576
rect 14558 40632 14624 40637
rect 14558 40576 14563 40632
rect 14619 40576 14624 40632
rect 14558 40571 14624 40576
rect 14858 40632 14924 40637
rect 14858 40576 14863 40632
rect 14919 40576 14924 40632
rect 14858 40571 14924 40576
rect 20300 40484 20500 40490
rect 21029 40484 21229 40489
rect 24034 40484 24234 40489
rect 20500 40286 21034 40484
rect 20300 40284 21034 40286
rect 21224 40284 24039 40484
rect 24229 40284 24234 40484
rect 20300 40280 20500 40284
rect 21029 40279 21229 40284
rect 24034 40279 24234 40284
rect 6500 40084 6700 40090
rect 13100 40084 13300 40090
rect 20900 40084 21100 40090
rect 21279 40084 21479 40089
rect 3720 40079 6500 40084
rect 3720 39889 3725 40079
rect 3915 39889 6021 40079
rect 6211 39889 6500 40079
rect 3720 39886 6500 39889
rect 6700 40079 13100 40084
rect 6700 39889 8141 40079
rect 8331 39889 10437 40079
rect 10627 39889 12557 40079
rect 12747 39889 13100 40079
rect 6700 39886 13100 39889
rect 13300 40079 15048 40084
rect 13300 39889 14853 40079
rect 15043 39889 15048 40079
rect 13300 39886 15048 39889
rect 3720 39884 15048 39886
rect 21100 39886 21284 40084
rect 20900 39884 21284 39886
rect 21474 39884 24139 40084
rect 6500 39880 6700 39884
rect 13100 39880 13300 39884
rect 20900 39880 21100 39884
rect 21279 39879 21479 39884
rect 7100 39684 7300 39690
rect 13700 39684 13900 39690
rect 3470 39679 7100 39684
rect 3470 39489 3475 39679
rect 3665 39489 6271 39679
rect 6461 39489 7100 39679
rect 3470 39486 7100 39489
rect 7300 39679 13700 39684
rect 7300 39489 7891 39679
rect 8081 39489 10687 39679
rect 10877 39489 12307 39679
rect 12497 39489 13700 39679
rect 7300 39486 13700 39489
rect 13900 39679 15298 39684
rect 13900 39489 15103 39679
rect 15293 39489 15298 39679
rect 13900 39486 15298 39489
rect 3470 39484 15298 39486
rect 7100 39480 7300 39484
rect 13700 39480 13900 39484
rect 20900 38484 21100 38490
rect 23784 38484 23984 38489
rect 21100 38286 23789 38484
rect 20900 38284 23789 38286
rect 23979 38284 24139 38484
rect 20900 38280 21100 38284
rect 23784 38279 23984 38284
rect 21633 37864 21699 37869
rect 21633 37808 21638 37864
rect 21694 37808 21699 37864
rect 21633 37803 21699 37808
rect 21933 37864 21999 37869
rect 21933 37808 21938 37864
rect 21994 37808 21999 37864
rect 21933 37803 21999 37808
rect 22233 37864 22299 37869
rect 22233 37808 22238 37864
rect 22294 37808 22299 37864
rect 22233 37803 22299 37808
rect 22533 37864 22599 37869
rect 22533 37808 22538 37864
rect 22594 37808 22599 37864
rect 22533 37803 22599 37808
rect 22833 37864 22899 37869
rect 22833 37808 22838 37864
rect 22894 37808 22899 37864
rect 22833 37803 22899 37808
rect 23133 37864 23199 37869
rect 23133 37808 23138 37864
rect 23194 37808 23199 37864
rect 23133 37803 23199 37808
rect 23433 37864 23499 37869
rect 23433 37808 23438 37864
rect 23494 37808 23499 37864
rect 23433 37803 23499 37808
rect 23733 37864 23799 37869
rect 23733 37808 23738 37864
rect 23794 37808 23799 37864
rect 23733 37803 23799 37808
rect 21636 37000 21696 37803
rect 21936 37200 21996 37803
rect 22236 37400 22296 37803
rect 22536 37400 22596 37803
rect 22236 37340 22377 37400
rect 21936 37140 22251 37200
rect 21636 36940 22125 37000
rect 22065 33280 22125 36940
rect 22191 33280 22251 37140
rect 22317 33280 22377 37340
rect 22443 37340 22596 37400
rect 22443 33280 22503 37340
rect 22836 37200 22896 37803
rect 22569 37140 22896 37200
rect 22569 33280 22629 37140
rect 23136 37000 23196 37803
rect 22695 36940 23196 37000
rect 22695 33280 22755 36940
rect 23436 36804 23496 37803
rect 22821 36744 23496 36804
rect 22821 33280 22881 36744
rect 23436 36740 23496 36744
rect 23736 36600 23796 37803
rect 22947 36540 23796 36600
rect 22947 33280 23007 36540
rect 7700 32127 7900 32133
rect 14300 32127 14500 32133
rect 20900 32127 21100 32133
rect 6065 31929 7700 32127
rect 7900 31929 14300 32127
rect 14500 31929 20900 32127
rect 21100 31929 21661 32127
rect 6065 31927 21661 31929
rect 7700 31923 7900 31927
rect 14300 31923 14500 31927
rect 20900 31923 21100 31927
rect 7100 31727 7300 31733
rect 13700 31727 13900 31733
rect 20300 31727 20500 31733
rect 6065 31529 7100 31727
rect 7300 31529 13700 31727
rect 13900 31529 20300 31727
rect 20500 31529 21661 31727
rect 6065 31527 21661 31529
rect 7100 31523 7300 31527
rect 13700 31523 13900 31527
rect 20300 31523 20500 31527
rect 6500 31327 6700 31333
rect 13100 31327 13300 31333
rect 19700 31327 19900 31333
rect 6065 31129 6500 31327
rect 6700 31129 13100 31327
rect 13300 31129 19700 31327
rect 19900 31129 21661 31327
rect 6065 31127 21661 31129
rect 6500 31123 6700 31127
rect 13100 31123 13300 31127
rect 19700 31123 19900 31127
rect 7700 27727 7900 27733
rect 14300 27727 14500 27733
rect 20900 27727 21100 27733
rect 6065 27529 7700 27727
rect 7900 27529 14300 27727
rect 14500 27529 20900 27727
rect 21100 27529 21661 27727
rect 6065 27527 21661 27529
rect 7700 27523 7900 27527
rect 14300 27523 14500 27527
rect 20900 27523 21100 27527
rect 7100 27327 7300 27333
rect 13700 27327 13900 27333
rect 20300 27327 20500 27333
rect 6065 27129 7100 27327
rect 7300 27129 13700 27327
rect 13900 27129 20300 27327
rect 20500 27129 21661 27327
rect 6065 27127 21661 27129
rect 7100 27123 7300 27127
rect 13700 27123 13900 27127
rect 20300 27123 20500 27127
rect 11899 26098 21682 26103
rect 11899 25928 21507 26098
rect 21677 25928 21682 26098
rect 11899 25923 21682 25928
rect 23012 26098 27414 26103
rect 23012 25928 23018 26098
rect 23188 25928 27414 26098
rect 23012 25923 27414 25928
rect 7700 18747 7900 18753
rect 14300 18747 14500 18753
rect 20900 18747 21100 18753
rect 6065 18549 7700 18747
rect 7900 18549 14300 18747
rect 14500 18549 20900 18747
rect 21100 18549 21661 18747
rect 6065 18547 21661 18549
rect 7700 18543 7900 18547
rect 14300 18543 14500 18547
rect 20900 18543 21100 18547
rect 7100 18347 7300 18353
rect 13700 18347 13900 18353
rect 20300 18347 20500 18353
rect 6065 18149 7100 18347
rect 7300 18149 13700 18347
rect 13900 18149 20300 18347
rect 20500 18149 21661 18347
rect 6065 18147 21661 18149
rect 7100 18143 7300 18147
rect 13700 18143 13900 18147
rect 20300 18143 20500 18147
rect 7700 12747 7900 12753
rect 14300 12747 14500 12753
rect 20900 12747 21100 12753
rect 6065 12549 7700 12747
rect 7900 12549 14300 12747
rect 14500 12549 20900 12747
rect 21100 12549 21661 12747
rect 6065 12547 21661 12549
rect 7700 12543 7900 12547
rect 14300 12543 14500 12547
rect 20900 12543 21100 12547
rect 7100 12347 7300 12353
rect 13700 12347 13900 12353
rect 20300 12347 20500 12353
rect 6065 12149 7100 12347
rect 7300 12149 13700 12347
rect 13900 12149 20300 12347
rect 20500 12149 21661 12347
rect 6065 12147 21661 12149
rect 7100 12143 7300 12147
rect 13700 12143 13900 12147
rect 20300 12143 20500 12147
rect 6500 11947 6700 11953
rect 13100 11947 13300 11953
rect 19700 11947 19900 11953
rect 6065 11749 6500 11947
rect 6700 11749 13100 11947
rect 13300 11749 19700 11947
rect 19900 11749 21661 11947
rect 6065 11747 21661 11749
rect 6500 11743 6700 11747
rect 13100 11743 13300 11747
rect 19700 11743 19900 11747
rect 27234 199 27414 25923
rect 27229 21 27235 199
rect 27413 21 27419 199
rect 27234 20 27414 21
<< via3 >>
rect 3004 44950 3068 45014
rect 3556 44950 3620 45014
rect 4108 44950 4172 45014
rect 4660 44950 4724 45014
rect 5212 44950 5276 45014
rect 5764 44950 5828 45014
rect 6316 44950 6380 45014
rect 6868 44950 6932 45014
rect 7420 44950 7484 45014
rect 7972 44950 8036 45014
rect 8524 44950 8588 45014
rect 9076 44950 9140 45014
rect 9628 44950 9692 45014
rect 10180 44950 10244 45014
rect 10732 44950 10796 45014
rect 11284 44950 11348 45014
rect 11836 44950 11900 45014
rect 12388 44950 12452 45014
rect 12940 44950 13004 45014
rect 13492 44950 13556 45014
rect 14044 44950 14108 45014
rect 14596 44950 14660 45014
rect 15148 44950 15212 45014
rect 15700 44950 15764 45014
rect 20668 44950 20732 45014
rect 21220 44950 21284 45014
rect 21772 44950 21836 45014
rect 22324 44950 22388 45014
rect 22876 44950 22940 45014
rect 23428 44950 23492 45014
rect 23980 44952 24044 45016
rect 24532 44950 24596 45014
rect 19700 40686 19900 40884
rect 20300 40286 20500 40484
rect 6500 39886 6700 40084
rect 13100 39886 13300 40084
rect 20900 39886 21100 40084
rect 7100 39486 7300 39684
rect 13700 39486 13900 39684
rect 20900 38286 21100 38484
rect 7700 31929 7900 32127
rect 14300 31929 14500 32127
rect 20900 31929 21100 32127
rect 7100 31529 7300 31727
rect 13700 31529 13900 31727
rect 20300 31529 20500 31727
rect 6500 31129 6700 31327
rect 13100 31129 13300 31327
rect 19700 31129 19900 31327
rect 7700 27529 7900 27727
rect 14300 27529 14500 27727
rect 20900 27529 21100 27727
rect 7100 27129 7300 27327
rect 13700 27129 13900 27327
rect 20300 27129 20500 27327
rect 7700 18549 7900 18747
rect 14300 18549 14500 18747
rect 20900 18549 21100 18747
rect 7100 18149 7300 18347
rect 13700 18149 13900 18347
rect 20300 18149 20500 18347
rect 7700 12549 7900 12747
rect 14300 12549 14500 12747
rect 20900 12549 21100 12747
rect 7100 12149 7300 12347
rect 13700 12149 13900 12347
rect 20300 12149 20500 12347
rect 6500 11749 6700 11947
rect 13100 11749 13300 11947
rect 19700 11749 19900 11947
rect 27235 21 27413 199
<< metal4 >>
rect 3006 45015 3066 45152
rect 3558 45015 3618 45152
rect 4110 45015 4170 45152
rect 4662 45015 4722 45152
rect 5214 45015 5274 45152
rect 5766 45015 5826 45152
rect 6318 45015 6378 45152
rect 6870 45015 6930 45152
rect 7422 45015 7482 45152
rect 7974 45015 8034 45152
rect 8526 45015 8586 45152
rect 9078 45015 9138 45152
rect 9630 45015 9690 45152
rect 10182 45015 10242 45152
rect 10734 45015 10794 45152
rect 11286 45015 11346 45152
rect 11838 45015 11898 45152
rect 12390 45015 12450 45152
rect 12942 45015 13002 45152
rect 13494 45015 13554 45152
rect 14046 45015 14106 45152
rect 14598 45015 14658 45152
rect 15150 45015 15210 45152
rect 15702 45015 15762 45152
rect 3003 45014 3069 45015
rect 3003 44950 3004 45014
rect 3068 44950 3069 45014
rect 3003 44949 3069 44950
rect 3555 45014 3621 45015
rect 3555 44950 3556 45014
rect 3620 44950 3621 45014
rect 3555 44949 3621 44950
rect 4107 45014 4173 45015
rect 4107 44950 4108 45014
rect 4172 44950 4173 45014
rect 4107 44949 4173 44950
rect 4659 45014 4725 45015
rect 4659 44950 4660 45014
rect 4724 44950 4725 45014
rect 4659 44949 4725 44950
rect 5211 45014 5277 45015
rect 5211 44950 5212 45014
rect 5276 44950 5277 45014
rect 5211 44949 5277 44950
rect 5763 45014 5829 45015
rect 5763 44950 5764 45014
rect 5828 44950 5829 45014
rect 5763 44949 5829 44950
rect 6315 45014 6381 45015
rect 6315 44950 6316 45014
rect 6380 44950 6381 45014
rect 6315 44949 6381 44950
rect 6867 45014 6933 45015
rect 6867 44950 6868 45014
rect 6932 44950 6933 45014
rect 6867 44949 6933 44950
rect 7419 45014 7485 45015
rect 7419 44950 7420 45014
rect 7484 44950 7485 45014
rect 7419 44949 7485 44950
rect 7971 45014 8037 45015
rect 7971 44950 7972 45014
rect 8036 44950 8037 45014
rect 7971 44949 8037 44950
rect 8523 45014 8589 45015
rect 8523 44950 8524 45014
rect 8588 44950 8589 45014
rect 8523 44949 8589 44950
rect 9075 45014 9141 45015
rect 9075 44950 9076 45014
rect 9140 44950 9141 45014
rect 9075 44949 9141 44950
rect 9627 45014 9693 45015
rect 9627 44950 9628 45014
rect 9692 44950 9693 45014
rect 9627 44949 9693 44950
rect 10179 45014 10245 45015
rect 10179 44950 10180 45014
rect 10244 44950 10245 45014
rect 10179 44949 10245 44950
rect 10731 45014 10797 45015
rect 10731 44950 10732 45014
rect 10796 44950 10797 45014
rect 10731 44949 10797 44950
rect 11283 45014 11349 45015
rect 11283 44950 11284 45014
rect 11348 44950 11349 45014
rect 11283 44949 11349 44950
rect 11835 45014 11901 45015
rect 11835 44950 11836 45014
rect 11900 44950 11901 45014
rect 11835 44949 11901 44950
rect 12387 45014 12453 45015
rect 12387 44950 12388 45014
rect 12452 44950 12453 45014
rect 12387 44949 12453 44950
rect 12939 45014 13005 45015
rect 12939 44950 12940 45014
rect 13004 44950 13005 45014
rect 12939 44949 13005 44950
rect 13491 45014 13557 45015
rect 13491 44950 13492 45014
rect 13556 44950 13557 45014
rect 13491 44949 13557 44950
rect 14043 45014 14109 45015
rect 14043 44950 14044 45014
rect 14108 44950 14109 45014
rect 14043 44949 14109 44950
rect 14595 45014 14661 45015
rect 14595 44950 14596 45014
rect 14660 44950 14661 45014
rect 14595 44949 14661 44950
rect 15147 45014 15213 45015
rect 15147 44950 15148 45014
rect 15212 44950 15213 45014
rect 15147 44949 15213 44950
rect 15699 45014 15765 45015
rect 15699 44950 15700 45014
rect 15764 44950 15765 45014
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 45015 20730 45152
rect 21222 45015 21282 45152
rect 21774 45015 21834 45152
rect 22326 45015 22386 45152
rect 22878 45015 22938 45152
rect 23430 45015 23490 45152
rect 23982 45017 24042 45152
rect 23979 45016 24045 45017
rect 20667 45014 20733 45015
rect 15699 44949 15765 44950
rect 20667 44950 20668 45014
rect 20732 44950 20733 45014
rect 20667 44949 20733 44950
rect 21219 45014 21285 45015
rect 21219 44950 21220 45014
rect 21284 44950 21285 45014
rect 21219 44949 21285 44950
rect 21771 45014 21837 45015
rect 21771 44950 21772 45014
rect 21836 44950 21837 45014
rect 21771 44949 21837 44950
rect 22323 45014 22389 45015
rect 22323 44950 22324 45014
rect 22388 44950 22389 45014
rect 22323 44949 22389 44950
rect 22875 45014 22941 45015
rect 22875 44950 22876 45014
rect 22940 44950 22941 45014
rect 22875 44949 22941 44950
rect 23427 45014 23493 45015
rect 23427 44950 23428 45014
rect 23492 44950 23493 45014
rect 23979 44952 23980 45016
rect 24044 44952 24045 45016
rect 24534 45015 24594 45152
rect 23979 44951 24045 44952
rect 24531 45014 24597 45015
rect 23427 44949 23493 44950
rect 24531 44950 24532 45014
rect 24596 44950 24597 45014
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 24531 44949 24597 44950
rect 6400 40084 6800 44152
rect 6400 39886 6500 40084
rect 6700 39886 6800 40084
rect 6400 31327 6800 39886
rect 6400 31129 6500 31327
rect 6700 31129 6800 31327
rect 6400 11947 6800 31129
rect 6400 11749 6500 11947
rect 6700 11749 6800 11947
rect 6400 1000 6800 11749
rect 7000 39684 7400 44152
rect 7000 39486 7100 39684
rect 7300 39486 7400 39684
rect 7000 31727 7400 39486
rect 7000 31529 7100 31727
rect 7300 31529 7400 31727
rect 7000 27327 7400 31529
rect 7000 27129 7100 27327
rect 7300 27129 7400 27327
rect 7000 18347 7400 27129
rect 7000 18149 7100 18347
rect 7300 18149 7400 18347
rect 7000 12347 7400 18149
rect 7000 12149 7100 12347
rect 7300 12149 7400 12347
rect 7000 1000 7400 12149
rect 7600 32127 8000 44152
rect 7600 31929 7700 32127
rect 7900 31929 8000 32127
rect 7600 27727 8000 31929
rect 7600 27529 7700 27727
rect 7900 27529 8000 27727
rect 7600 18747 8000 27529
rect 7600 18549 7700 18747
rect 7900 18549 8000 18747
rect 7600 12747 8000 18549
rect 7600 12549 7700 12747
rect 7900 12549 8000 12747
rect 7600 1000 8000 12549
rect 13000 40084 13400 44152
rect 13000 39886 13100 40084
rect 13300 39886 13400 40084
rect 13000 31327 13400 39886
rect 13000 31129 13100 31327
rect 13300 31129 13400 31327
rect 13000 11947 13400 31129
rect 13000 11749 13100 11947
rect 13300 11749 13400 11947
rect 13000 1000 13400 11749
rect 13600 39684 14000 44152
rect 13600 39486 13700 39684
rect 13900 39486 14000 39684
rect 13600 31727 14000 39486
rect 13600 31529 13700 31727
rect 13900 31529 14000 31727
rect 13600 27327 14000 31529
rect 13600 27129 13700 27327
rect 13900 27129 14000 27327
rect 13600 18347 14000 27129
rect 13600 18149 13700 18347
rect 13900 18149 14000 18347
rect 13600 12347 14000 18149
rect 13600 12149 13700 12347
rect 13900 12149 14000 12347
rect 13600 1000 14000 12149
rect 14200 32127 14600 44152
rect 14200 31929 14300 32127
rect 14500 31929 14600 32127
rect 14200 27727 14600 31929
rect 14200 27529 14300 27727
rect 14500 27529 14600 27727
rect 14200 18747 14600 27529
rect 14200 18549 14300 18747
rect 14500 18549 14600 18747
rect 14200 12747 14600 18549
rect 14200 12549 14300 12747
rect 14500 12549 14600 12747
rect 14200 1000 14600 12549
rect 19600 40884 20000 44152
rect 19600 40686 19700 40884
rect 19900 40686 20000 40884
rect 19600 31327 20000 40686
rect 19600 31129 19700 31327
rect 19900 31129 20000 31327
rect 19600 11947 20000 31129
rect 19600 11749 19700 11947
rect 19900 11749 20000 11947
rect 19600 1000 20000 11749
rect 20200 40484 20600 44152
rect 20200 40286 20300 40484
rect 20500 40286 20600 40484
rect 20200 31727 20600 40286
rect 20200 31529 20300 31727
rect 20500 31529 20600 31727
rect 20200 27327 20600 31529
rect 20200 27129 20300 27327
rect 20500 27129 20600 27327
rect 20200 18347 20600 27129
rect 20200 18149 20300 18347
rect 20500 18149 20600 18347
rect 20200 12347 20600 18149
rect 20200 12149 20300 12347
rect 20500 12149 20600 12347
rect 20200 1000 20600 12149
rect 20800 40084 21200 44152
rect 20800 39886 20900 40084
rect 21100 39886 21200 40084
rect 20800 38484 21200 39886
rect 20800 38286 20900 38484
rect 21100 38286 21200 38484
rect 20800 32127 21200 38286
rect 20800 31929 20900 32127
rect 21100 31929 21200 32127
rect 20800 27727 21200 31929
rect 20800 27529 20900 27727
rect 21100 27529 21200 27727
rect 20800 18747 21200 27529
rect 20800 18549 20900 18747
rect 21100 18549 21200 18747
rect 20800 12747 21200 18549
rect 20800 12549 20900 12747
rect 21100 12549 21200 12747
rect 20800 1000 21200 12549
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 199 27414 200
rect 27234 21 27235 199
rect 27413 21 27414 199
rect 27234 0 27414 21
use dac  dac_0
timestamp 1748333863
transform 1 0 6065 0 1 12147
box -4 -396 16945 21433
use shifters  shifters_0
timestamp 1748318706
transform 1 0 21337 0 1 37600
box -213 0 2802 3976
use tie_lows  tie_lows_0
timestamp 1748318706
transform 1 0 12462 0 1 40284
box -110 0 2786 1292
use tie_lows  tie_lows_1
timestamp 1748318706
transform 1 0 8046 0 1 40284
box -110 0 2786 1292
use tie_lows  tie_lows_2
timestamp 1748318706
transform 1 0 3630 0 1 40284
box -110 0 2786 1292
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 6400 1000 6800 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 7000 1000 7400 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 7600 1000 8000 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 19600 1000 20000 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 20200 1000 20600 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 20800 1000 21200 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 13000 1000 13400 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 13600 1000 14000 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 14200 1000 14600 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
