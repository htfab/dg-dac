magic
tech sky130A
magscale 1 2
timestamp 1748076069
<< metal1 >>
rect 148 5744 15448 5802
rect 972 4785 1006 5629
rect 1872 4785 1906 5629
rect 2772 4785 2806 5629
rect 3672 4785 3706 5629
rect 4572 4785 4606 5629
rect 5472 4785 5506 5629
rect 6372 4785 6406 5629
rect 7272 4785 7306 5629
rect 8172 4785 8206 5629
rect 9072 4785 9106 5629
rect 9972 4785 10006 5629
rect 10872 4785 10906 5629
rect 11772 4785 11806 5629
rect 12672 4785 12706 5629
rect 13572 4785 13606 5629
rect 14472 4785 14506 5629
rect 15372 4785 15406 5629
rect 272 4760 324 4766
rect 272 4702 324 4708
rect 572 4760 624 4766
rect 572 4702 624 4708
rect 1172 4760 1224 4766
rect 1172 4702 1224 4708
rect 1472 4760 1524 4766
rect 1472 4702 1524 4708
rect 2072 4760 2124 4766
rect 2072 4702 2124 4708
rect 2372 4760 2424 4766
rect 2372 4702 2424 4708
rect 2972 4760 3024 4766
rect 2972 4702 3024 4708
rect 3272 4760 3324 4766
rect 3272 4702 3324 4708
rect 3872 4760 3924 4766
rect 3872 4702 3924 4708
rect 4172 4760 4224 4766
rect 4172 4702 4224 4708
rect 4772 4760 4824 4766
rect 4772 4702 4824 4708
rect 5072 4760 5124 4766
rect 5072 4702 5124 4708
rect 5672 4760 5724 4766
rect 5672 4702 5724 4708
rect 5972 4760 6024 4766
rect 5972 4702 6024 4708
rect 6572 4760 6624 4766
rect 6572 4702 6624 4708
rect 6872 4760 6924 4766
rect 6872 4702 6924 4708
rect 7472 4760 7524 4766
rect 7472 4702 7524 4708
rect 7772 4760 7824 4766
rect 7772 4702 7824 4708
rect 8372 4760 8424 4766
rect 8372 4702 8424 4708
rect 8672 4760 8724 4766
rect 8672 4702 8724 4708
rect 9272 4760 9324 4766
rect 9272 4702 9324 4708
rect 9572 4760 9624 4766
rect 9572 4702 9624 4708
rect 10172 4760 10224 4766
rect 10172 4702 10224 4708
rect 10472 4760 10524 4766
rect 10472 4702 10524 4708
rect 11072 4760 11124 4766
rect 11072 4702 11124 4708
rect 11372 4760 11424 4766
rect 11372 4702 11424 4708
rect 11972 4760 12024 4766
rect 11972 4702 12024 4708
rect 12272 4760 12324 4766
rect 12272 4702 12324 4708
rect 12872 4760 12924 4766
rect 12872 4702 12924 4708
rect 13172 4760 13224 4766
rect 13172 4702 13224 4708
rect 13772 4760 13824 4766
rect 13772 4702 13824 4708
rect 14072 4760 14124 4766
rect 14072 4702 14124 4708
rect 14672 4760 14724 4766
rect 14672 4702 14724 4708
rect 14972 4760 15024 4766
rect 14972 4702 15024 4708
rect 272 4670 324 4673
rect 14972 4670 15024 4673
rect 148 4667 15448 4670
rect 148 4615 272 4667
rect 324 4615 14972 4667
rect 15024 4615 15448 4667
rect 148 4612 15448 4615
rect 272 4609 324 4612
rect 14972 4609 15024 4612
rect 572 4542 624 4548
rect 1172 4542 1224 4548
rect 624 4499 1172 4533
rect 572 4484 624 4490
rect 1172 4484 1224 4490
rect 1472 4465 1524 4471
rect 2072 4465 2124 4471
rect 1524 4422 2072 4456
rect 1472 4407 1524 4413
rect 2072 4407 2124 4413
rect 2372 4388 2424 4394
rect 2972 4388 3024 4394
rect 2424 4345 2972 4379
rect 2372 4330 2424 4336
rect 2972 4330 3024 4336
rect 3272 4311 3324 4317
rect 3872 4311 3924 4317
rect 3324 4268 3872 4302
rect 3272 4253 3324 4259
rect 3872 4253 3924 4259
rect 4172 4234 4224 4240
rect 4772 4234 4824 4240
rect 4224 4191 4772 4225
rect 4172 4176 4224 4182
rect 4772 4176 4824 4182
rect 5072 4157 5124 4163
rect 5672 4157 5724 4163
rect 5124 4114 5672 4148
rect 5072 4099 5124 4105
rect 5672 4099 5724 4105
rect 5972 4080 6024 4086
rect 6572 4080 6624 4086
rect 6024 4037 6572 4071
rect 5972 4022 6024 4028
rect 6572 4022 6624 4028
rect 6872 4003 6924 4009
rect 7472 4003 7524 4009
rect 6924 3960 7472 3994
rect 6872 3945 6924 3951
rect 7472 3945 7524 3951
rect 7772 3926 7824 3932
rect 8372 3926 8424 3932
rect 7824 3883 8372 3917
rect 7772 3868 7824 3874
rect 8372 3868 8424 3874
rect 8672 3849 8724 3855
rect 9272 3849 9324 3855
rect 8724 3806 9272 3840
rect 8672 3791 8724 3797
rect 9272 3791 9324 3797
rect 9572 3772 9624 3778
rect 10172 3772 10224 3778
rect 9624 3729 10172 3763
rect 9572 3714 9624 3720
rect 10172 3714 10224 3720
rect 10472 3695 10524 3701
rect 11072 3695 11124 3701
rect 10524 3652 11072 3686
rect 10472 3637 10524 3643
rect 11072 3637 11124 3643
rect 11372 3618 11424 3624
rect 11972 3618 12024 3624
rect 11424 3575 11972 3609
rect 11372 3560 11424 3566
rect 11972 3560 12024 3566
rect 12272 3541 12324 3547
rect 12872 3541 12924 3547
rect 12324 3498 12872 3532
rect 12272 3483 12324 3489
rect 12872 3483 12924 3489
rect 13172 3464 13224 3470
rect 13772 3464 13824 3470
rect 13224 3421 13772 3455
rect 13172 3406 13224 3412
rect 13772 3406 13824 3412
rect 14072 3387 14124 3393
rect 14672 3387 14724 3393
rect 14124 3344 14672 3378
rect 14072 3329 14124 3335
rect 14672 3329 14724 3335
<< via1 >>
rect 272 4708 324 4760
rect 572 4708 624 4760
rect 1172 4708 1224 4760
rect 1472 4708 1524 4760
rect 2072 4708 2124 4760
rect 2372 4708 2424 4760
rect 2972 4708 3024 4760
rect 3272 4708 3324 4760
rect 3872 4708 3924 4760
rect 4172 4708 4224 4760
rect 4772 4708 4824 4760
rect 5072 4708 5124 4760
rect 5672 4708 5724 4760
rect 5972 4708 6024 4760
rect 6572 4708 6624 4760
rect 6872 4708 6924 4760
rect 7472 4708 7524 4760
rect 7772 4708 7824 4760
rect 8372 4708 8424 4760
rect 8672 4708 8724 4760
rect 9272 4708 9324 4760
rect 9572 4708 9624 4760
rect 10172 4708 10224 4760
rect 10472 4708 10524 4760
rect 11072 4708 11124 4760
rect 11372 4708 11424 4760
rect 11972 4708 12024 4760
rect 12272 4708 12324 4760
rect 12872 4708 12924 4760
rect 13172 4708 13224 4760
rect 13772 4708 13824 4760
rect 14072 4708 14124 4760
rect 14672 4708 14724 4760
rect 14972 4708 15024 4760
rect 272 4615 324 4667
rect 14972 4615 15024 4667
rect 572 4490 624 4542
rect 1172 4490 1224 4542
rect 1472 4413 1524 4465
rect 2072 4413 2124 4465
rect 2372 4336 2424 4388
rect 2972 4336 3024 4388
rect 3272 4259 3324 4311
rect 3872 4259 3924 4311
rect 4172 4182 4224 4234
rect 4772 4182 4824 4234
rect 5072 4105 5124 4157
rect 5672 4105 5724 4157
rect 5972 4028 6024 4080
rect 6572 4028 6624 4080
rect 6872 3951 6924 4003
rect 7472 3951 7524 4003
rect 7772 3874 7824 3926
rect 8372 3874 8424 3926
rect 8672 3797 8724 3849
rect 9272 3797 9324 3849
rect 9572 3720 9624 3772
rect 10172 3720 10224 3772
rect 10472 3643 10524 3695
rect 11072 3643 11124 3695
rect 11372 3566 11424 3618
rect 11972 3566 12024 3618
rect 12272 3489 12324 3541
rect 12872 3489 12924 3541
rect 13172 3412 13224 3464
rect 13772 3412 13824 3464
rect 14072 3335 14124 3387
rect 14672 3335 14724 3387
<< metal2 >>
rect 266 4708 272 4760
rect 324 4708 330 4760
rect 566 4708 572 4760
rect 624 4708 630 4760
rect 1166 4708 1172 4760
rect 1224 4708 1230 4760
rect 1466 4708 1472 4760
rect 1524 4708 1530 4760
rect 2066 4708 2072 4760
rect 2124 4708 2130 4760
rect 2366 4708 2372 4760
rect 2424 4708 2430 4760
rect 2966 4708 2972 4760
rect 3024 4708 3030 4760
rect 3266 4708 3272 4760
rect 3324 4708 3330 4760
rect 3866 4708 3872 4760
rect 3924 4708 3930 4760
rect 4166 4708 4172 4760
rect 4224 4708 4230 4760
rect 4766 4708 4772 4760
rect 4824 4708 4830 4760
rect 5066 4708 5072 4760
rect 5124 4708 5130 4760
rect 5666 4708 5672 4760
rect 5724 4708 5730 4760
rect 5966 4708 5972 4760
rect 6024 4708 6030 4760
rect 6566 4708 6572 4760
rect 6624 4708 6630 4760
rect 6866 4708 6872 4760
rect 6924 4708 6930 4760
rect 7466 4708 7472 4760
rect 7524 4708 7530 4760
rect 7766 4708 7772 4760
rect 7824 4708 7830 4760
rect 8366 4708 8372 4760
rect 8424 4708 8430 4760
rect 8666 4708 8672 4760
rect 8724 4708 8730 4760
rect 9266 4708 9272 4760
rect 9324 4708 9330 4760
rect 9566 4708 9572 4760
rect 9624 4708 9630 4760
rect 10166 4708 10172 4760
rect 10224 4708 10230 4760
rect 10466 4708 10472 4760
rect 10524 4708 10530 4760
rect 11066 4708 11072 4760
rect 11124 4708 11130 4760
rect 11366 4708 11372 4760
rect 11424 4708 11430 4760
rect 11966 4708 11972 4760
rect 12024 4708 12030 4760
rect 12266 4708 12272 4760
rect 12324 4708 12330 4760
rect 12866 4708 12872 4760
rect 12924 4708 12930 4760
rect 13166 4708 13172 4760
rect 13224 4708 13230 4760
rect 13766 4708 13772 4760
rect 13824 4708 13830 4760
rect 14066 4708 14072 4760
rect 14124 4708 14130 4760
rect 14666 4708 14672 4760
rect 14724 4708 14730 4760
rect 14966 4708 14972 4760
rect 15024 4708 15030 4760
rect 281 4667 315 4708
rect 266 4615 272 4667
rect 324 4615 330 4667
rect 581 4542 615 4708
rect 1181 4542 1215 4708
rect 566 4490 572 4542
rect 624 4490 630 4542
rect 1166 4490 1172 4542
rect 1224 4490 1230 4542
rect 1481 4465 1515 4708
rect 2081 4465 2115 4708
rect 1466 4413 1472 4465
rect 1524 4413 1530 4465
rect 2066 4413 2072 4465
rect 2124 4413 2130 4465
rect 2381 4388 2415 4708
rect 2981 4388 3015 4708
rect 2366 4336 2372 4388
rect 2424 4336 2430 4388
rect 2966 4336 2972 4388
rect 3024 4336 3030 4388
rect 3281 4311 3315 4708
rect 3881 4311 3915 4708
rect 3266 4259 3272 4311
rect 3324 4259 3330 4311
rect 3866 4259 3872 4311
rect 3924 4259 3930 4311
rect 4181 4234 4215 4708
rect 4781 4234 4815 4708
rect 4166 4182 4172 4234
rect 4224 4182 4230 4234
rect 4766 4182 4772 4234
rect 4824 4182 4830 4234
rect 5081 4157 5115 4708
rect 5681 4157 5715 4708
rect 5066 4105 5072 4157
rect 5124 4105 5130 4157
rect 5666 4105 5672 4157
rect 5724 4105 5730 4157
rect 5981 4080 6015 4708
rect 6581 4080 6615 4708
rect 5966 4028 5972 4080
rect 6024 4028 6030 4080
rect 6566 4028 6572 4080
rect 6624 4028 6630 4080
rect 6881 4003 6915 4708
rect 7481 4003 7515 4708
rect 6866 3951 6872 4003
rect 6924 3951 6930 4003
rect 7466 3951 7472 4003
rect 7524 3951 7530 4003
rect 7781 3926 7815 4708
rect 8381 3926 8415 4708
rect 7766 3874 7772 3926
rect 7824 3874 7830 3926
rect 8366 3874 8372 3926
rect 8424 3874 8430 3926
rect 8681 3849 8715 4708
rect 9281 3849 9315 4708
rect 8666 3797 8672 3849
rect 8724 3797 8730 3849
rect 9266 3797 9272 3849
rect 9324 3797 9330 3849
rect 9581 3772 9615 4708
rect 10181 3772 10215 4708
rect 9566 3720 9572 3772
rect 9624 3720 9630 3772
rect 10166 3720 10172 3772
rect 10224 3720 10230 3772
rect 10481 3695 10515 4708
rect 11081 3695 11115 4708
rect 10466 3643 10472 3695
rect 10524 3643 10530 3695
rect 11066 3643 11072 3695
rect 11124 3643 11130 3695
rect 11381 3618 11415 4708
rect 11981 3618 12015 4708
rect 11366 3566 11372 3618
rect 11424 3566 11430 3618
rect 11966 3566 11972 3618
rect 12024 3566 12030 3618
rect 12281 3541 12315 4708
rect 12881 3541 12915 4708
rect 12266 3489 12272 3541
rect 12324 3489 12330 3541
rect 12866 3489 12872 3541
rect 12924 3489 12930 3541
rect 13181 3464 13215 4708
rect 13781 3464 13815 4708
rect 13166 3412 13172 3464
rect 13224 3412 13230 3464
rect 13766 3412 13772 3464
rect 13824 3412 13830 3464
rect 14081 3387 14115 4708
rect 14681 3387 14715 4708
rect 14981 4667 15015 4708
rect 14966 4615 14972 4667
rect 15024 4615 15030 4667
rect 14066 3335 14072 3387
rect 14124 3335 14130 3387
rect 14666 3335 14672 3387
rect 14724 3335 14730 3387
use multi_or2  multi_or2_0
timestamp 1748065934
transform 1 0 0 0 1 4576
box 0 0 15596 1292
<< labels >>
flabel metal1 972 4785 1006 5629 1 FreeSans 128 0 0 0 C[0]
port 18 nsew signal output
flabel metal1 1872 4785 1906 5629 1 FreeSans 128 0 0 0 C[1]
port 19 nsew signal output
flabel metal1 2772 4785 2806 5629 1 FreeSans 128 0 0 0 C[2]
port 20 nsew signal output
flabel metal1 3672 4785 3706 5629 1 FreeSans 128 0 0 0 C[3]
port 21 nsew signal output
flabel metal1 4572 4785 4606 5629 1 FreeSans 128 0 0 0 C[4]
port 22 nsew signal output
flabel metal1 5472 4785 5506 5629 1 FreeSans 128 0 0 0 C[5]
port 23 nsew signal output
flabel metal1 6372 4785 6406 5629 1 FreeSans 128 0 0 0 C[6]
port 24 nsew signal output
flabel metal1 7272 4785 7306 5629 1 FreeSans 128 0 0 0 C[7]
port 25 nsew signal output
flabel metal1 8172 4785 8206 5629 1 FreeSans 128 0 0 0 C[8]
port 26 nsew signal output
flabel metal1 9072 4785 9106 5629 1 FreeSans 128 0 0 0 C[9]
port 27 nsew signal output
flabel metal1 9972 4785 10006 5629 1 FreeSans 128 0 0 0 C[10]
port 28 nsew signal output
flabel metal1 10872 4785 10906 5629 1 FreeSans 128 0 0 0 C[11]
port 29 nsew signal output
flabel metal1 11772 4785 11806 5629 1 FreeSans 128 0 0 0 C[12]
port 30 nsew signal output
flabel metal1 12672 4785 12706 5629 1 FreeSans 128 0 0 0 C[13]
port 31 nsew signal output
flabel metal1 13572 4785 13606 5629 1 FreeSans 128 0 0 0 C[14]
port 32 nsew signal output
flabel metal1 14472 4785 14506 5629 1 FreeSans 128 0 0 0 C[15]
port 33 nsew signal output
flabel metal1 15372 4785 15406 5629 1 FreeSans 128 0 0 0 C[16]
port 34 nsew signal output
flabel metal1 148 4612 15448 4670 0 FreeSans 256 0 0 0 VSS
port 0 nsew ground bidirectional
flabel metal1 148 5744 15448 5802 0 FreeSans 256 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal1 624 4499 1172 4533 0 FreeSans 256 0 0 0 U[0]
port 2 nsew signal input
flabel metal1 1524 4422 2072 4456 0 FreeSans 256 0 0 0 U[1]
port 3 nsew signal input
flabel metal1 2424 4345 2972 4379 0 FreeSans 256 0 0 0 U[2]
port 4 nsew signal input
flabel metal1 3324 4268 3872 4302 0 FreeSans 256 0 0 0 U[3]
port 5 nsew signal input
flabel metal1 4224 4191 4772 4225 0 FreeSans 256 0 0 0 U[4]
port 6 nsew signal input
flabel metal1 5124 4114 5672 4148 0 FreeSans 256 0 0 0 U[5]
port 7 nsew signal input
flabel metal1 6024 4037 6572 4071 0 FreeSans 256 0 0 0 U[6]
port 8 nsew signal input
flabel metal1 6924 3960 7472 3994 0 FreeSans 256 0 0 0 U[7]
port 9 nsew signal input
flabel metal1 7824 3883 8372 3917 0 FreeSans 256 0 0 0 U[8]
port 10 nsew signal input
flabel metal1 8724 3806 9272 3840 0 FreeSans 256 0 0 0 U[9]
port 11 nsew signal input
flabel metal1 9624 3729 10172 3763 0 FreeSans 256 0 0 0 U[10]
port 12 nsew signal input
flabel metal1 10524 3652 11072 3686 0 FreeSans 256 0 0 0 U[11]
port 13 nsew signal input
flabel metal1 11424 3575 11972 3609 0 FreeSans 256 0 0 0 U[12]
port 14 nsew signal input
flabel metal1 12324 3498 12872 3532 0 FreeSans 256 0 0 0 U[13]
port 15 nsew signal input
flabel metal1 13224 3421 13772 3455 0 FreeSans 256 0 0 0 U[14]
port 16 nsew signal input
flabel metal1 14124 3344 14672 3378 0 FreeSans 256 0 0 0 U[15]
port 17 nsew signal input
<< end >>
