magic
tech sky130A
magscale 1 2
timestamp 1748299483
<< metal1 >>
rect 148 1168 2524 1226
rect 281 898 315 1130
rect 266 846 272 898
rect 324 846 330 898
rect 281 141 315 846
rect 581 714 615 1130
rect 866 846 872 898
rect 924 846 930 898
rect 1257 846 1263 898
rect 1315 846 1321 898
rect 2066 846 2072 898
rect 2124 846 2130 898
rect 566 662 572 714
rect 624 662 630 714
rect 1166 662 1172 714
rect 1224 662 1230 714
rect 1857 662 1863 714
rect 1915 662 1921 714
rect 2366 662 2372 714
rect 2424 662 2430 714
rect 357 478 363 530
rect 415 478 421 530
rect 581 141 615 662
rect 1466 478 1472 530
rect 1524 478 1530 530
rect 657 294 663 346
rect 715 294 721 346
rect 1766 294 1772 346
rect 1824 294 1830 346
rect 2472 209 2506 1053
rect 148 36 2524 94
<< via1 >>
rect 272 846 324 898
rect 872 846 924 898
rect 1263 846 1315 898
rect 2072 846 2124 898
rect 572 662 624 714
rect 1172 662 1224 714
rect 1863 662 1915 714
rect 2372 662 2424 714
rect 363 478 415 530
rect 1472 478 1524 530
rect 663 294 715 346
rect 1772 294 1824 346
<< metal2 >>
rect 272 898 324 904
rect 872 898 924 904
rect 324 855 872 889
rect 272 840 324 846
rect 872 840 924 846
rect 1263 898 1315 904
rect 2072 898 2124 904
rect 1315 855 2072 889
rect 1263 840 1315 846
rect 2072 840 2124 846
rect 572 714 624 720
rect 1172 714 1224 720
rect 624 671 1172 705
rect 572 656 624 662
rect 1172 656 1224 662
rect 1863 714 1915 720
rect 2372 714 2424 720
rect 1915 671 2372 705
rect 1863 656 1915 662
rect 2372 656 2424 662
rect 363 530 415 536
rect 1472 530 1524 536
rect 415 487 1472 521
rect 363 472 415 478
rect 1472 472 1524 478
rect 663 346 715 352
rect 1772 346 1824 352
rect 715 303 1772 337
rect 663 288 715 294
rect 1772 288 1824 294
use inverter_raw  inverter_raw_0
timestamp 1748299149
transform 1 0 60 0 1 0
box 88 36 388 1226
use inverter_raw  inverter_raw_1
timestamp 1748299149
transform 1 0 360 0 1 0
box 88 36 388 1226
use nor2_raw  nor2_raw_0
timestamp 1748299149
transform 1 0 660 0 1 0
box 88 36 664 1226
use nor2_raw  nor2_raw_1
timestamp 1748299149
transform 1 0 1260 0 1 0
box 88 36 664 1226
use nor2_raw  nor2_raw_2
timestamp 1748299149
transform 1 0 1860 0 1 0
box 88 36 664 1226
<< labels >>
flabel metal1 281 141 315 1130 0 FreeSans 256 0 0 0 A
port 2 nsew signal input
flabel metal1 581 141 615 1130 0 FreeSans 256 0 0 0 B
port 3 nsew signal input
flabel metal1 2472 209 2506 1053 0 FreeSans 128 0 0 0 OUT
port 4 nsew signal output
flabel metal1 148 36 2524 94 0 FreeSans 256 0 0 0 VSS
port 0 nsew ground bidirectional
flabel metal1 148 1168 2524 1226 0 FreeSans 256 0 0 0 VDD
port 1 nsew power bidirectional
<< end >>
