magic
tech sky130A
magscale 1 2
timestamp 1748060222
<< locali >>
rect -63 3414 37 3420
rect -63 3356 -51 3414
rect 25 3402 37 3414
rect 2552 3414 2652 3420
rect 2552 3402 2564 3414
rect 25 3368 124 3402
rect 2452 3368 2564 3402
rect 25 3356 37 3368
rect -63 3350 37 3356
rect 2552 3356 2564 3368
rect 2640 3356 2652 3414
rect 2552 3350 2652 3356
rect -63 3204 37 3210
rect -63 3146 -51 3204
rect 25 3192 37 3204
rect 2552 3204 2652 3210
rect 2552 3192 2564 3204
rect 25 3158 124 3192
rect 2452 3158 2564 3192
rect 25 3146 37 3158
rect -63 3140 37 3146
rect 2552 3146 2564 3158
rect 2640 3146 2652 3204
rect 2552 3140 2652 3146
rect -63 2072 37 2078
rect -63 2014 -51 2072
rect 25 2060 37 2072
rect 2552 2072 2652 2078
rect 2552 2060 2564 2072
rect 25 2026 124 2060
rect 2452 2026 2564 2060
rect 25 2014 37 2026
rect -63 2008 37 2014
rect 2552 2014 2564 2026
rect 2640 2014 2652 2072
rect 2552 2008 2652 2014
rect -63 1862 37 1868
rect -63 1804 -51 1862
rect 25 1850 37 1862
rect 2552 1862 2652 1868
rect 2552 1850 2564 1862
rect 25 1816 124 1850
rect 2452 1816 2564 1850
rect 25 1804 37 1816
rect -63 1798 37 1804
rect 2552 1804 2564 1816
rect 2640 1804 2652 1862
rect 2552 1798 2652 1804
rect -63 730 37 736
rect -63 672 -51 730
rect 25 718 37 730
rect 2552 730 2652 736
rect 2552 718 2564 730
rect 25 684 124 718
rect 2452 684 2564 718
rect 25 672 37 684
rect -63 666 37 672
rect 2552 672 2564 684
rect 2640 672 2652 730
rect 2552 666 2652 672
rect -63 520 37 526
rect -63 462 -51 520
rect 25 508 37 520
rect 2552 520 2652 526
rect 2552 508 2564 520
rect 25 474 124 508
rect 2452 474 2564 508
rect 25 462 37 474
rect -63 456 37 462
rect 2552 462 2564 474
rect 2640 462 2652 520
rect 2552 456 2652 462
<< viali >>
rect -51 3356 25 3414
rect 2564 3356 2640 3414
rect -51 3146 25 3204
rect 2564 3146 2640 3204
rect -51 2014 25 2072
rect 2564 2014 2640 2072
rect -51 1804 25 1862
rect 2564 1804 2640 1862
rect -51 672 25 730
rect 2564 672 2640 730
rect -51 462 25 520
rect 2564 462 2640 520
<< metal1 >>
rect -63 3910 37 3916
rect 2552 3910 2652 3916
rect -63 3852 -51 3910
rect 25 3852 2564 3910
rect 2640 3852 2652 3910
rect -63 3846 37 3852
rect 2552 3846 2652 3852
rect -63 3414 37 3420
rect -63 3356 -51 3414
rect 25 3356 37 3414
rect -63 3350 37 3356
rect -213 3204 37 3210
rect -213 3146 -201 3204
rect -125 3146 -51 3204
rect 25 3146 37 3204
rect -213 3140 37 3146
rect 221 2819 255 3820
rect 521 2819 555 3820
rect 821 2819 855 3820
rect 1121 2819 1155 3820
rect 1421 2819 1455 3820
rect 1721 2819 1755 3820
rect 2021 2819 2055 3820
rect 2321 2819 2355 3820
rect 2552 3414 2652 3420
rect 2552 3356 2564 3414
rect 2640 3356 2652 3414
rect 2552 3350 2652 3356
rect 2552 3204 2802 3210
rect 2552 3146 2564 3204
rect 2640 3146 2714 3204
rect 2790 3146 2802 3204
rect 2552 3140 2802 3146
rect -213 2778 -113 2784
rect 2702 2778 2802 2784
rect -213 2720 -201 2778
rect -125 2720 2714 2778
rect 2790 2720 2802 2778
rect -213 2714 -113 2720
rect 2702 2714 2802 2720
rect -63 2568 37 2574
rect 2552 2568 2652 2574
rect -63 2510 -51 2568
rect 25 2510 2564 2568
rect 2640 2510 2652 2568
rect -63 2504 37 2510
rect 2552 2504 2652 2510
rect -63 2072 37 2078
rect -63 2014 -51 2072
rect 25 2014 37 2072
rect -63 2008 37 2014
rect 2552 2072 2652 2078
rect 2552 2014 2564 2072
rect 2640 2014 2652 2072
rect 2552 2008 2652 2014
rect -213 1862 37 1868
rect -213 1804 -201 1862
rect -125 1804 -51 1862
rect 25 1804 37 1862
rect -213 1798 37 1804
rect 2552 1862 2802 1868
rect 2552 1804 2564 1862
rect 2640 1804 2714 1862
rect 2790 1804 2802 1862
rect 2552 1798 2802 1804
rect -213 1436 -113 1442
rect 2702 1436 2802 1442
rect -213 1378 -201 1436
rect -125 1378 2714 1436
rect 2790 1378 2802 1436
rect -213 1372 -113 1378
rect 2702 1372 2802 1378
rect -63 1226 37 1232
rect 2552 1226 2652 1232
rect -63 1168 -51 1226
rect 25 1168 2564 1226
rect 2640 1168 2652 1226
rect -63 1162 37 1168
rect 2552 1162 2652 1168
rect -63 730 37 736
rect -63 672 -51 730
rect 25 672 37 730
rect -63 666 37 672
rect -213 520 37 526
rect -213 462 -201 520
rect -125 462 -51 520
rect 25 462 37 520
rect -213 456 37 462
rect 312 209 346 1053
rect 612 209 646 1053
rect 912 209 946 1053
rect 1212 209 1246 1053
rect 1512 209 1546 1053
rect 1812 209 1846 1053
rect 2112 209 2146 1053
rect 2412 209 2446 1053
rect 2552 730 2652 736
rect 2552 672 2564 730
rect 2640 672 2652 730
rect 2552 666 2652 672
rect 2552 520 2802 526
rect 2552 462 2564 520
rect 2640 462 2714 520
rect 2790 462 2802 520
rect 2552 456 2802 462
rect -213 94 -113 100
rect 2702 94 2802 100
rect -213 36 -201 94
rect -125 36 2714 94
rect 2790 36 2802 94
rect -213 30 -113 36
rect 2702 30 2802 36
<< via1 >>
rect -51 3852 25 3910
rect 2564 3852 2640 3910
rect -51 3356 25 3414
rect -201 3146 -125 3204
rect 2564 3356 2640 3414
rect 2714 3146 2790 3204
rect -201 2720 -125 2778
rect 2714 2720 2790 2778
rect -51 2510 25 2568
rect 2564 2510 2640 2568
rect -51 2014 25 2072
rect 2564 2014 2640 2072
rect -201 1804 -125 1862
rect 2714 1804 2790 1862
rect -201 1378 -125 1436
rect 2714 1378 2790 1436
rect -51 1168 25 1226
rect 2564 1168 2640 1226
rect -51 672 25 730
rect -201 462 -125 520
rect 2564 672 2640 730
rect 2714 462 2790 520
rect -201 36 -125 94
rect 2714 36 2790 94
<< metal2 >>
rect -213 3204 -113 3976
rect -213 3146 -201 3204
rect -125 3146 -113 3204
rect -213 2778 -113 3146
rect -213 2720 -201 2778
rect -125 2720 -113 2778
rect -63 3910 37 3976
rect -63 3852 -51 3910
rect 25 3852 37 3910
rect -63 3414 37 3852
rect -63 3356 -51 3414
rect 25 3356 37 3414
rect -63 2721 37 3356
rect 2552 3910 2652 3976
rect 2552 3852 2564 3910
rect 2640 3852 2652 3910
rect 2552 3414 2652 3852
rect 2552 3356 2564 3414
rect 2640 3356 2652 3414
rect 2552 2721 2652 3356
rect 2702 3204 2802 3976
rect 2702 3146 2714 3204
rect 2790 3146 2802 3204
rect 2702 2778 2802 3146
rect -213 1862 -113 2720
rect 2702 2720 2714 2778
rect 2790 2720 2802 2778
rect -213 1804 -201 1862
rect -125 1804 -113 1862
rect -213 1436 -113 1804
rect -213 1378 -201 1436
rect -125 1378 -113 1436
rect -213 520 -113 1378
rect -213 462 -201 520
rect -125 462 -113 520
rect -213 94 -113 462
rect -213 36 -201 94
rect -125 36 -113 94
rect -213 0 -113 36
rect -63 2568 37 2574
rect -63 2510 -51 2568
rect 25 2510 37 2568
rect -63 2072 37 2510
rect -63 2014 -51 2072
rect 25 2014 37 2072
rect -63 1226 37 2014
rect -63 1168 -51 1226
rect 25 1168 37 1226
rect -63 730 37 1168
rect -63 672 -51 730
rect 25 672 37 730
rect -63 0 37 672
rect 2552 2568 2652 2574
rect 2552 2510 2564 2568
rect 2640 2510 2652 2568
rect 2552 2072 2652 2510
rect 2552 2014 2564 2072
rect 2640 2014 2652 2072
rect 2552 1226 2652 2014
rect 2552 1168 2564 1226
rect 2640 1168 2652 1226
rect 2552 730 2652 1168
rect 2552 672 2564 730
rect 2640 672 2652 730
rect 2552 0 2652 672
rect 2702 1862 2802 2720
rect 2702 1804 2714 1862
rect 2790 1804 2802 1862
rect 2702 1436 2802 1804
rect 2702 1378 2714 1436
rect 2790 1378 2802 1436
rect 2702 520 2802 1378
rect 2702 462 2714 520
rect 2790 462 2802 520
rect 2702 94 2802 462
rect 2702 36 2714 94
rect 2790 36 2802 94
rect 2702 0 2802 36
use shifter_raw  shifter_raw_1
array 0 7 300 0 0 6127
timestamp 1748060222
transform 1 0 0 0 1 0
box 88 36 388 3910
use transistor_pair_bus_8  transistor_pair_bus_8_0
timestamp 1740627177
transform 1 0 0 0 1 0
box -60 0 2636 1292
use transistor_pair_bus_8  transistor_pair_bus_8_1
timestamp 1740627177
transform 1 0 0 0 1 1342
box -60 0 2636 1292
use transistor_pair_bus_8  transistor_pair_bus_8_2
timestamp 1740627177
transform 1 0 0 0 1 2684
box -60 0 2636 1292
<< labels >>
flabel metal1 2321 2819 2355 3820 1 FreeSans 400 0 0 0 IN[0]
port 1 n signal default
flabel metal1 2021 2819 2055 3820 1 FreeSans 400 0 0 0 IN[1]
port 2 n signal default
flabel metal1 1721 2819 1755 3820 1 FreeSans 400 0 0 0 IN[2]
port 3 n signal default
flabel metal1 1421 2819 1455 3820 1 FreeSans 400 0 0 0 IN[3]
port 4 n signal default
flabel metal1 1121 2819 1155 3820 1 FreeSans 400 0 0 0 IN[4]
port 5 n signal default
flabel metal1 821 2819 855 3820 1 FreeSans 400 0 0 0 IN[5]
port 6 n signal default
flabel metal1 521 2819 555 3820 1 FreeSans 400 0 0 0 IN[6]
port 7 n signal default
flabel metal1 221 2819 255 3820 1 FreeSans 400 0 0 0 IN[7]
port 8 n signal default
flabel metal1 2412 209 2446 1053 1 FreeSans 400 0 0 0 OUT[0]
port 9 n signal default
flabel metal1 2112 209 2146 1053 1 FreeSans 400 0 0 0 OUT[1]
port 10 n signal default
flabel metal1 1812 209 1846 1053 1 FreeSans 400 0 0 0 OUT[2]
port 11 n signal default
flabel metal1 1512 209 1546 1053 1 FreeSans 400 0 0 0 OUT[3]
port 12 n signal default
flabel metal1 1212 209 1246 1053 1 FreeSans 400 0 0 0 OUT[4]
port 13 n signal default
flabel metal1 912 209 946 1053 1 FreeSans 400 0 0 0 OUT[5]
port 14 n signal default
flabel metal1 612 209 646 1053 1 FreeSans 400 0 0 0 OUT[6]
port 15 n signal default
flabel metal1 312 209 346 1053 1 FreeSans 400 0 0 0 OUT[7]
port 16 n signal default
flabel metal2 -213 0 -113 3976 1 FreeSans 400 0 0 0 VSS
port 17 n ground bidirectional
flabel metal2 -63 2721 37 3976 1 FreeSans 400 0 0 0 IVDD
port 18 n power bidirectional
flabel metal2 -63 0 37 2568 1 FreeSans 400 0 0 0 OVDD
port 19 n power bidirectional
<< end >>
