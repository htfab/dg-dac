magic
tech sky130A
magscale 1 2
timestamp 1748309517
<< nwell >>
rect 0 954 5540 2076
<< pwell >>
rect 10 0 5540 904
<< mvnmos >>
rect 236 561 336 691
rect 512 561 612 691
rect 788 561 888 691
rect 1064 561 1164 691
rect 1340 561 1440 691
rect 1616 561 1716 691
rect 1892 561 1992 691
rect 2168 561 2268 691
rect 2444 561 2544 691
rect 2720 561 2820 691
rect 2996 561 3096 691
rect 3272 561 3372 691
rect 3548 561 3648 691
rect 3824 561 3924 691
rect 4100 561 4200 691
rect 4376 561 4476 691
rect 4652 561 4752 691
rect 4928 561 5028 691
rect 5204 561 5304 691
rect 236 213 336 343
rect 512 213 612 343
rect 788 213 888 343
rect 1064 213 1164 343
rect 1340 213 1440 343
rect 1616 213 1716 343
rect 1892 213 1992 343
rect 2168 213 2268 343
rect 2444 213 2544 343
rect 2720 213 2820 343
rect 2996 213 3096 343
rect 3272 213 3372 343
rect 3548 213 3648 343
rect 3824 213 3924 343
rect 4100 213 4200 343
rect 4376 213 4476 343
rect 4652 213 4752 343
rect 4928 213 5028 343
rect 5204 213 5304 343
<< mvpmos >>
rect 236 1633 336 1833
rect 512 1633 612 1833
rect 788 1633 888 1833
rect 1064 1633 1164 1833
rect 1340 1633 1440 1833
rect 1616 1633 1716 1833
rect 1892 1633 1992 1833
rect 2168 1633 2268 1833
rect 2444 1633 2544 1833
rect 2720 1633 2820 1833
rect 2996 1633 3096 1833
rect 3272 1633 3372 1833
rect 3548 1633 3648 1833
rect 3824 1633 3924 1833
rect 4100 1633 4200 1833
rect 4376 1633 4476 1833
rect 4652 1633 4752 1833
rect 4928 1633 5028 1833
rect 5204 1633 5304 1833
rect 236 1197 336 1397
rect 512 1197 612 1397
rect 788 1197 888 1397
rect 1064 1197 1164 1397
rect 1340 1197 1440 1397
rect 1616 1197 1716 1397
rect 1892 1197 1992 1397
rect 2168 1197 2268 1397
rect 2444 1197 2544 1397
rect 2720 1197 2820 1397
rect 2996 1197 3096 1397
rect 3272 1197 3372 1397
rect 3548 1197 3648 1397
rect 3824 1197 3924 1397
rect 4100 1197 4200 1397
rect 4376 1197 4476 1397
rect 4652 1197 4752 1397
rect 4928 1197 5028 1397
rect 5204 1197 5304 1397
<< mvndiff >>
rect 178 679 236 691
rect 178 573 190 679
rect 224 573 236 679
rect 178 561 236 573
rect 336 679 394 691
rect 336 573 348 679
rect 382 573 394 679
rect 336 561 394 573
rect 454 679 512 691
rect 454 573 466 679
rect 500 573 512 679
rect 454 561 512 573
rect 612 679 670 691
rect 612 573 624 679
rect 658 573 670 679
rect 612 561 670 573
rect 730 679 788 691
rect 730 573 742 679
rect 776 573 788 679
rect 730 561 788 573
rect 888 679 946 691
rect 888 573 900 679
rect 934 573 946 679
rect 888 561 946 573
rect 1006 679 1064 691
rect 1006 573 1018 679
rect 1052 573 1064 679
rect 1006 561 1064 573
rect 1164 679 1222 691
rect 1164 573 1176 679
rect 1210 573 1222 679
rect 1164 561 1222 573
rect 1282 679 1340 691
rect 1282 573 1294 679
rect 1328 573 1340 679
rect 1282 561 1340 573
rect 1440 679 1498 691
rect 1440 573 1452 679
rect 1486 573 1498 679
rect 1440 561 1498 573
rect 1558 679 1616 691
rect 1558 573 1570 679
rect 1604 573 1616 679
rect 1558 561 1616 573
rect 1716 679 1774 691
rect 1716 573 1728 679
rect 1762 573 1774 679
rect 1716 561 1774 573
rect 1834 679 1892 691
rect 1834 573 1846 679
rect 1880 573 1892 679
rect 1834 561 1892 573
rect 1992 679 2050 691
rect 1992 573 2004 679
rect 2038 573 2050 679
rect 1992 561 2050 573
rect 2110 679 2168 691
rect 2110 573 2122 679
rect 2156 573 2168 679
rect 2110 561 2168 573
rect 2268 679 2326 691
rect 2268 573 2280 679
rect 2314 573 2326 679
rect 2268 561 2326 573
rect 2386 679 2444 691
rect 2386 573 2398 679
rect 2432 573 2444 679
rect 2386 561 2444 573
rect 2544 679 2602 691
rect 2544 573 2556 679
rect 2590 573 2602 679
rect 2544 561 2602 573
rect 2662 679 2720 691
rect 2662 573 2674 679
rect 2708 573 2720 679
rect 2662 561 2720 573
rect 2820 679 2878 691
rect 2820 573 2832 679
rect 2866 573 2878 679
rect 2820 561 2878 573
rect 2938 679 2996 691
rect 2938 573 2950 679
rect 2984 573 2996 679
rect 2938 561 2996 573
rect 3096 679 3154 691
rect 3096 573 3108 679
rect 3142 573 3154 679
rect 3096 561 3154 573
rect 3214 679 3272 691
rect 3214 573 3226 679
rect 3260 573 3272 679
rect 3214 561 3272 573
rect 3372 679 3430 691
rect 3372 573 3384 679
rect 3418 573 3430 679
rect 3372 561 3430 573
rect 3490 679 3548 691
rect 3490 573 3502 679
rect 3536 573 3548 679
rect 3490 561 3548 573
rect 3648 679 3706 691
rect 3648 573 3660 679
rect 3694 573 3706 679
rect 3648 561 3706 573
rect 3766 679 3824 691
rect 3766 573 3778 679
rect 3812 573 3824 679
rect 3766 561 3824 573
rect 3924 679 3982 691
rect 3924 573 3936 679
rect 3970 573 3982 679
rect 3924 561 3982 573
rect 4042 679 4100 691
rect 4042 573 4054 679
rect 4088 573 4100 679
rect 4042 561 4100 573
rect 4200 679 4258 691
rect 4200 573 4212 679
rect 4246 573 4258 679
rect 4200 561 4258 573
rect 4318 679 4376 691
rect 4318 573 4330 679
rect 4364 573 4376 679
rect 4318 561 4376 573
rect 4476 679 4534 691
rect 4476 573 4488 679
rect 4522 573 4534 679
rect 4476 561 4534 573
rect 4594 679 4652 691
rect 4594 573 4606 679
rect 4640 573 4652 679
rect 4594 561 4652 573
rect 4752 679 4810 691
rect 4752 573 4764 679
rect 4798 573 4810 679
rect 4752 561 4810 573
rect 4870 679 4928 691
rect 4870 573 4882 679
rect 4916 573 4928 679
rect 4870 561 4928 573
rect 5028 679 5086 691
rect 5028 573 5040 679
rect 5074 573 5086 679
rect 5028 561 5086 573
rect 5146 679 5204 691
rect 5146 573 5158 679
rect 5192 573 5204 679
rect 5146 561 5204 573
rect 5304 679 5362 691
rect 5304 573 5316 679
rect 5350 573 5362 679
rect 5304 561 5362 573
rect 178 331 236 343
rect 178 225 190 331
rect 224 225 236 331
rect 178 213 236 225
rect 336 331 394 343
rect 336 225 348 331
rect 382 225 394 331
rect 336 213 394 225
rect 454 331 512 343
rect 454 225 466 331
rect 500 225 512 331
rect 454 213 512 225
rect 612 331 670 343
rect 612 225 624 331
rect 658 225 670 331
rect 612 213 670 225
rect 730 331 788 343
rect 730 225 742 331
rect 776 225 788 331
rect 730 213 788 225
rect 888 331 946 343
rect 888 225 900 331
rect 934 225 946 331
rect 888 213 946 225
rect 1006 331 1064 343
rect 1006 225 1018 331
rect 1052 225 1064 331
rect 1006 213 1064 225
rect 1164 331 1222 343
rect 1164 225 1176 331
rect 1210 225 1222 331
rect 1164 213 1222 225
rect 1282 331 1340 343
rect 1282 225 1294 331
rect 1328 225 1340 331
rect 1282 213 1340 225
rect 1440 331 1498 343
rect 1440 225 1452 331
rect 1486 225 1498 331
rect 1440 213 1498 225
rect 1558 331 1616 343
rect 1558 225 1570 331
rect 1604 225 1616 331
rect 1558 213 1616 225
rect 1716 331 1774 343
rect 1716 225 1728 331
rect 1762 225 1774 331
rect 1716 213 1774 225
rect 1834 331 1892 343
rect 1834 225 1846 331
rect 1880 225 1892 331
rect 1834 213 1892 225
rect 1992 331 2050 343
rect 1992 225 2004 331
rect 2038 225 2050 331
rect 1992 213 2050 225
rect 2110 331 2168 343
rect 2110 225 2122 331
rect 2156 225 2168 331
rect 2110 213 2168 225
rect 2268 331 2326 343
rect 2268 225 2280 331
rect 2314 225 2326 331
rect 2268 213 2326 225
rect 2386 331 2444 343
rect 2386 225 2398 331
rect 2432 225 2444 331
rect 2386 213 2444 225
rect 2544 331 2602 343
rect 2544 225 2556 331
rect 2590 225 2602 331
rect 2544 213 2602 225
rect 2662 331 2720 343
rect 2662 225 2674 331
rect 2708 225 2720 331
rect 2662 213 2720 225
rect 2820 331 2878 343
rect 2820 225 2832 331
rect 2866 225 2878 331
rect 2820 213 2878 225
rect 2938 331 2996 343
rect 2938 225 2950 331
rect 2984 225 2996 331
rect 2938 213 2996 225
rect 3096 331 3154 343
rect 3096 225 3108 331
rect 3142 225 3154 331
rect 3096 213 3154 225
rect 3214 331 3272 343
rect 3214 225 3226 331
rect 3260 225 3272 331
rect 3214 213 3272 225
rect 3372 331 3430 343
rect 3372 225 3384 331
rect 3418 225 3430 331
rect 3372 213 3430 225
rect 3490 331 3548 343
rect 3490 225 3502 331
rect 3536 225 3548 331
rect 3490 213 3548 225
rect 3648 331 3706 343
rect 3648 225 3660 331
rect 3694 225 3706 331
rect 3648 213 3706 225
rect 3766 331 3824 343
rect 3766 225 3778 331
rect 3812 225 3824 331
rect 3766 213 3824 225
rect 3924 331 3982 343
rect 3924 225 3936 331
rect 3970 225 3982 331
rect 3924 213 3982 225
rect 4042 331 4100 343
rect 4042 225 4054 331
rect 4088 225 4100 331
rect 4042 213 4100 225
rect 4200 331 4258 343
rect 4200 225 4212 331
rect 4246 225 4258 331
rect 4200 213 4258 225
rect 4318 331 4376 343
rect 4318 225 4330 331
rect 4364 225 4376 331
rect 4318 213 4376 225
rect 4476 331 4534 343
rect 4476 225 4488 331
rect 4522 225 4534 331
rect 4476 213 4534 225
rect 4594 331 4652 343
rect 4594 225 4606 331
rect 4640 225 4652 331
rect 4594 213 4652 225
rect 4752 331 4810 343
rect 4752 225 4764 331
rect 4798 225 4810 331
rect 4752 213 4810 225
rect 4870 331 4928 343
rect 4870 225 4882 331
rect 4916 225 4928 331
rect 4870 213 4928 225
rect 5028 331 5086 343
rect 5028 225 5040 331
rect 5074 225 5086 331
rect 5028 213 5086 225
rect 5146 331 5204 343
rect 5146 225 5158 331
rect 5192 225 5204 331
rect 5146 213 5204 225
rect 5304 331 5362 343
rect 5304 225 5316 331
rect 5350 225 5362 331
rect 5304 213 5362 225
<< mvpdiff >>
rect 178 1821 236 1833
rect 178 1645 190 1821
rect 224 1645 236 1821
rect 178 1633 236 1645
rect 336 1821 394 1833
rect 336 1645 348 1821
rect 382 1645 394 1821
rect 336 1633 394 1645
rect 454 1821 512 1833
rect 454 1645 466 1821
rect 500 1645 512 1821
rect 454 1633 512 1645
rect 612 1821 670 1833
rect 612 1645 624 1821
rect 658 1645 670 1821
rect 612 1633 670 1645
rect 730 1821 788 1833
rect 730 1645 742 1821
rect 776 1645 788 1821
rect 730 1633 788 1645
rect 888 1821 946 1833
rect 888 1645 900 1821
rect 934 1645 946 1821
rect 888 1633 946 1645
rect 1006 1821 1064 1833
rect 1006 1645 1018 1821
rect 1052 1645 1064 1821
rect 1006 1633 1064 1645
rect 1164 1821 1222 1833
rect 1164 1645 1176 1821
rect 1210 1645 1222 1821
rect 1164 1633 1222 1645
rect 1282 1821 1340 1833
rect 1282 1645 1294 1821
rect 1328 1645 1340 1821
rect 1282 1633 1340 1645
rect 1440 1821 1498 1833
rect 1440 1645 1452 1821
rect 1486 1645 1498 1821
rect 1440 1633 1498 1645
rect 1558 1821 1616 1833
rect 1558 1645 1570 1821
rect 1604 1645 1616 1821
rect 1558 1633 1616 1645
rect 1716 1821 1774 1833
rect 1716 1645 1728 1821
rect 1762 1645 1774 1821
rect 1716 1633 1774 1645
rect 1834 1821 1892 1833
rect 1834 1645 1846 1821
rect 1880 1645 1892 1821
rect 1834 1633 1892 1645
rect 1992 1821 2050 1833
rect 1992 1645 2004 1821
rect 2038 1645 2050 1821
rect 1992 1633 2050 1645
rect 2110 1821 2168 1833
rect 2110 1645 2122 1821
rect 2156 1645 2168 1821
rect 2110 1633 2168 1645
rect 2268 1821 2326 1833
rect 2268 1645 2280 1821
rect 2314 1645 2326 1821
rect 2268 1633 2326 1645
rect 2386 1821 2444 1833
rect 2386 1645 2398 1821
rect 2432 1645 2444 1821
rect 2386 1633 2444 1645
rect 2544 1821 2602 1833
rect 2544 1645 2556 1821
rect 2590 1645 2602 1821
rect 2544 1633 2602 1645
rect 2662 1821 2720 1833
rect 2662 1645 2674 1821
rect 2708 1645 2720 1821
rect 2662 1633 2720 1645
rect 2820 1821 2878 1833
rect 2820 1645 2832 1821
rect 2866 1645 2878 1821
rect 2820 1633 2878 1645
rect 2938 1821 2996 1833
rect 2938 1645 2950 1821
rect 2984 1645 2996 1821
rect 2938 1633 2996 1645
rect 3096 1821 3154 1833
rect 3096 1645 3108 1821
rect 3142 1645 3154 1821
rect 3096 1633 3154 1645
rect 3214 1821 3272 1833
rect 3214 1645 3226 1821
rect 3260 1645 3272 1821
rect 3214 1633 3272 1645
rect 3372 1821 3430 1833
rect 3372 1645 3384 1821
rect 3418 1645 3430 1821
rect 3372 1633 3430 1645
rect 3490 1821 3548 1833
rect 3490 1645 3502 1821
rect 3536 1645 3548 1821
rect 3490 1633 3548 1645
rect 3648 1821 3706 1833
rect 3648 1645 3660 1821
rect 3694 1645 3706 1821
rect 3648 1633 3706 1645
rect 3766 1821 3824 1833
rect 3766 1645 3778 1821
rect 3812 1645 3824 1821
rect 3766 1633 3824 1645
rect 3924 1821 3982 1833
rect 3924 1645 3936 1821
rect 3970 1645 3982 1821
rect 3924 1633 3982 1645
rect 4042 1821 4100 1833
rect 4042 1645 4054 1821
rect 4088 1645 4100 1821
rect 4042 1633 4100 1645
rect 4200 1821 4258 1833
rect 4200 1645 4212 1821
rect 4246 1645 4258 1821
rect 4200 1633 4258 1645
rect 4318 1821 4376 1833
rect 4318 1645 4330 1821
rect 4364 1645 4376 1821
rect 4318 1633 4376 1645
rect 4476 1821 4534 1833
rect 4476 1645 4488 1821
rect 4522 1645 4534 1821
rect 4476 1633 4534 1645
rect 4594 1821 4652 1833
rect 4594 1645 4606 1821
rect 4640 1645 4652 1821
rect 4594 1633 4652 1645
rect 4752 1821 4810 1833
rect 4752 1645 4764 1821
rect 4798 1645 4810 1821
rect 4752 1633 4810 1645
rect 4870 1821 4928 1833
rect 4870 1645 4882 1821
rect 4916 1645 4928 1821
rect 4870 1633 4928 1645
rect 5028 1821 5086 1833
rect 5028 1645 5040 1821
rect 5074 1645 5086 1821
rect 5028 1633 5086 1645
rect 5146 1821 5204 1833
rect 5146 1645 5158 1821
rect 5192 1645 5204 1821
rect 5146 1633 5204 1645
rect 5304 1821 5362 1833
rect 5304 1645 5316 1821
rect 5350 1645 5362 1821
rect 5304 1633 5362 1645
rect 178 1385 236 1397
rect 178 1209 190 1385
rect 224 1209 236 1385
rect 178 1197 236 1209
rect 336 1385 394 1397
rect 336 1209 348 1385
rect 382 1209 394 1385
rect 336 1197 394 1209
rect 454 1385 512 1397
rect 454 1209 466 1385
rect 500 1209 512 1385
rect 454 1197 512 1209
rect 612 1385 670 1397
rect 612 1209 624 1385
rect 658 1209 670 1385
rect 612 1197 670 1209
rect 730 1385 788 1397
rect 730 1209 742 1385
rect 776 1209 788 1385
rect 730 1197 788 1209
rect 888 1385 946 1397
rect 888 1209 900 1385
rect 934 1209 946 1385
rect 888 1197 946 1209
rect 1006 1385 1064 1397
rect 1006 1209 1018 1385
rect 1052 1209 1064 1385
rect 1006 1197 1064 1209
rect 1164 1385 1222 1397
rect 1164 1209 1176 1385
rect 1210 1209 1222 1385
rect 1164 1197 1222 1209
rect 1282 1385 1340 1397
rect 1282 1209 1294 1385
rect 1328 1209 1340 1385
rect 1282 1197 1340 1209
rect 1440 1385 1498 1397
rect 1440 1209 1452 1385
rect 1486 1209 1498 1385
rect 1440 1197 1498 1209
rect 1558 1385 1616 1397
rect 1558 1209 1570 1385
rect 1604 1209 1616 1385
rect 1558 1197 1616 1209
rect 1716 1385 1774 1397
rect 1716 1209 1728 1385
rect 1762 1209 1774 1385
rect 1716 1197 1774 1209
rect 1834 1385 1892 1397
rect 1834 1209 1846 1385
rect 1880 1209 1892 1385
rect 1834 1197 1892 1209
rect 1992 1385 2050 1397
rect 1992 1209 2004 1385
rect 2038 1209 2050 1385
rect 1992 1197 2050 1209
rect 2110 1385 2168 1397
rect 2110 1209 2122 1385
rect 2156 1209 2168 1385
rect 2110 1197 2168 1209
rect 2268 1385 2326 1397
rect 2268 1209 2280 1385
rect 2314 1209 2326 1385
rect 2268 1197 2326 1209
rect 2386 1385 2444 1397
rect 2386 1209 2398 1385
rect 2432 1209 2444 1385
rect 2386 1197 2444 1209
rect 2544 1385 2602 1397
rect 2544 1209 2556 1385
rect 2590 1209 2602 1385
rect 2544 1197 2602 1209
rect 2662 1385 2720 1397
rect 2662 1209 2674 1385
rect 2708 1209 2720 1385
rect 2662 1197 2720 1209
rect 2820 1385 2878 1397
rect 2820 1209 2832 1385
rect 2866 1209 2878 1385
rect 2820 1197 2878 1209
rect 2938 1385 2996 1397
rect 2938 1209 2950 1385
rect 2984 1209 2996 1385
rect 2938 1197 2996 1209
rect 3096 1385 3154 1397
rect 3096 1209 3108 1385
rect 3142 1209 3154 1385
rect 3096 1197 3154 1209
rect 3214 1385 3272 1397
rect 3214 1209 3226 1385
rect 3260 1209 3272 1385
rect 3214 1197 3272 1209
rect 3372 1385 3430 1397
rect 3372 1209 3384 1385
rect 3418 1209 3430 1385
rect 3372 1197 3430 1209
rect 3490 1385 3548 1397
rect 3490 1209 3502 1385
rect 3536 1209 3548 1385
rect 3490 1197 3548 1209
rect 3648 1385 3706 1397
rect 3648 1209 3660 1385
rect 3694 1209 3706 1385
rect 3648 1197 3706 1209
rect 3766 1385 3824 1397
rect 3766 1209 3778 1385
rect 3812 1209 3824 1385
rect 3766 1197 3824 1209
rect 3924 1385 3982 1397
rect 3924 1209 3936 1385
rect 3970 1209 3982 1385
rect 3924 1197 3982 1209
rect 4042 1385 4100 1397
rect 4042 1209 4054 1385
rect 4088 1209 4100 1385
rect 4042 1197 4100 1209
rect 4200 1385 4258 1397
rect 4200 1209 4212 1385
rect 4246 1209 4258 1385
rect 4200 1197 4258 1209
rect 4318 1385 4376 1397
rect 4318 1209 4330 1385
rect 4364 1209 4376 1385
rect 4318 1197 4376 1209
rect 4476 1385 4534 1397
rect 4476 1209 4488 1385
rect 4522 1209 4534 1385
rect 4476 1197 4534 1209
rect 4594 1385 4652 1397
rect 4594 1209 4606 1385
rect 4640 1209 4652 1385
rect 4594 1197 4652 1209
rect 4752 1385 4810 1397
rect 4752 1209 4764 1385
rect 4798 1209 4810 1385
rect 4752 1197 4810 1209
rect 4870 1385 4928 1397
rect 4870 1209 4882 1385
rect 4916 1209 4928 1385
rect 4870 1197 4928 1209
rect 5028 1385 5086 1397
rect 5028 1209 5040 1385
rect 5074 1209 5086 1385
rect 5028 1197 5086 1209
rect 5146 1385 5204 1397
rect 5146 1209 5158 1385
rect 5192 1209 5204 1385
rect 5146 1197 5204 1209
rect 5304 1385 5362 1397
rect 5304 1209 5316 1385
rect 5350 1209 5362 1385
rect 5304 1197 5362 1209
<< mvndiffc >>
rect 190 573 224 679
rect 348 573 382 679
rect 466 573 500 679
rect 624 573 658 679
rect 742 573 776 679
rect 900 573 934 679
rect 1018 573 1052 679
rect 1176 573 1210 679
rect 1294 573 1328 679
rect 1452 573 1486 679
rect 1570 573 1604 679
rect 1728 573 1762 679
rect 1846 573 1880 679
rect 2004 573 2038 679
rect 2122 573 2156 679
rect 2280 573 2314 679
rect 2398 573 2432 679
rect 2556 573 2590 679
rect 2674 573 2708 679
rect 2832 573 2866 679
rect 2950 573 2984 679
rect 3108 573 3142 679
rect 3226 573 3260 679
rect 3384 573 3418 679
rect 3502 573 3536 679
rect 3660 573 3694 679
rect 3778 573 3812 679
rect 3936 573 3970 679
rect 4054 573 4088 679
rect 4212 573 4246 679
rect 4330 573 4364 679
rect 4488 573 4522 679
rect 4606 573 4640 679
rect 4764 573 4798 679
rect 4882 573 4916 679
rect 5040 573 5074 679
rect 5158 573 5192 679
rect 5316 573 5350 679
rect 190 225 224 331
rect 348 225 382 331
rect 466 225 500 331
rect 624 225 658 331
rect 742 225 776 331
rect 900 225 934 331
rect 1018 225 1052 331
rect 1176 225 1210 331
rect 1294 225 1328 331
rect 1452 225 1486 331
rect 1570 225 1604 331
rect 1728 225 1762 331
rect 1846 225 1880 331
rect 2004 225 2038 331
rect 2122 225 2156 331
rect 2280 225 2314 331
rect 2398 225 2432 331
rect 2556 225 2590 331
rect 2674 225 2708 331
rect 2832 225 2866 331
rect 2950 225 2984 331
rect 3108 225 3142 331
rect 3226 225 3260 331
rect 3384 225 3418 331
rect 3502 225 3536 331
rect 3660 225 3694 331
rect 3778 225 3812 331
rect 3936 225 3970 331
rect 4054 225 4088 331
rect 4212 225 4246 331
rect 4330 225 4364 331
rect 4488 225 4522 331
rect 4606 225 4640 331
rect 4764 225 4798 331
rect 4882 225 4916 331
rect 5040 225 5074 331
rect 5158 225 5192 331
rect 5316 225 5350 331
<< mvpdiffc >>
rect 190 1645 224 1821
rect 348 1645 382 1821
rect 466 1645 500 1821
rect 624 1645 658 1821
rect 742 1645 776 1821
rect 900 1645 934 1821
rect 1018 1645 1052 1821
rect 1176 1645 1210 1821
rect 1294 1645 1328 1821
rect 1452 1645 1486 1821
rect 1570 1645 1604 1821
rect 1728 1645 1762 1821
rect 1846 1645 1880 1821
rect 2004 1645 2038 1821
rect 2122 1645 2156 1821
rect 2280 1645 2314 1821
rect 2398 1645 2432 1821
rect 2556 1645 2590 1821
rect 2674 1645 2708 1821
rect 2832 1645 2866 1821
rect 2950 1645 2984 1821
rect 3108 1645 3142 1821
rect 3226 1645 3260 1821
rect 3384 1645 3418 1821
rect 3502 1645 3536 1821
rect 3660 1645 3694 1821
rect 3778 1645 3812 1821
rect 3936 1645 3970 1821
rect 4054 1645 4088 1821
rect 4212 1645 4246 1821
rect 4330 1645 4364 1821
rect 4488 1645 4522 1821
rect 4606 1645 4640 1821
rect 4764 1645 4798 1821
rect 4882 1645 4916 1821
rect 5040 1645 5074 1821
rect 5158 1645 5192 1821
rect 5316 1645 5350 1821
rect 190 1209 224 1385
rect 348 1209 382 1385
rect 466 1209 500 1385
rect 624 1209 658 1385
rect 742 1209 776 1385
rect 900 1209 934 1385
rect 1018 1209 1052 1385
rect 1176 1209 1210 1385
rect 1294 1209 1328 1385
rect 1452 1209 1486 1385
rect 1570 1209 1604 1385
rect 1728 1209 1762 1385
rect 1846 1209 1880 1385
rect 2004 1209 2038 1385
rect 2122 1209 2156 1385
rect 2280 1209 2314 1385
rect 2398 1209 2432 1385
rect 2556 1209 2590 1385
rect 2674 1209 2708 1385
rect 2832 1209 2866 1385
rect 2950 1209 2984 1385
rect 3108 1209 3142 1385
rect 3226 1209 3260 1385
rect 3384 1209 3418 1385
rect 3502 1209 3536 1385
rect 3660 1209 3694 1385
rect 3778 1209 3812 1385
rect 3936 1209 3970 1385
rect 4054 1209 4088 1385
rect 4212 1209 4246 1385
rect 4330 1209 4364 1385
rect 4488 1209 4522 1385
rect 4606 1209 4640 1385
rect 4764 1209 4798 1385
rect 4882 1209 4916 1385
rect 5040 1209 5074 1385
rect 5158 1209 5192 1385
rect 5316 1209 5350 1385
<< mvpsubdiff >>
rect 46 856 5504 868
rect 46 822 172 856
rect 400 822 448 856
rect 676 822 724 856
rect 952 822 1000 856
rect 1228 822 1276 856
rect 1504 822 1552 856
rect 1780 822 1828 856
rect 2056 822 2104 856
rect 2332 822 2380 856
rect 2608 822 2656 856
rect 2884 822 2932 856
rect 3160 822 3208 856
rect 3436 822 3484 856
rect 3712 822 3760 856
rect 3988 822 4036 856
rect 4264 822 4312 856
rect 4540 822 4588 856
rect 4816 822 4864 856
rect 5092 822 5140 856
rect 5368 822 5504 856
rect 46 810 5504 822
rect 46 760 104 810
rect 46 144 58 760
rect 92 144 104 760
rect 5446 760 5504 810
rect 46 94 104 144
rect 5446 144 5458 760
rect 5492 144 5504 760
rect 5446 94 5504 144
rect 46 82 5504 94
rect 46 48 172 82
rect 400 48 448 82
rect 676 48 724 82
rect 952 48 1000 82
rect 1228 48 1276 82
rect 1504 48 1552 82
rect 1780 48 1828 82
rect 2056 48 2104 82
rect 2332 48 2380 82
rect 2608 48 2656 82
rect 2884 48 2932 82
rect 3160 48 3208 82
rect 3436 48 3484 82
rect 3712 48 3760 82
rect 3988 48 4036 82
rect 4264 48 4312 82
rect 4540 48 4588 82
rect 4816 48 4864 82
rect 5092 48 5140 82
rect 5368 48 5504 82
rect 46 36 5504 48
<< mvnsubdiff >>
rect 66 1998 5474 2010
rect 66 1964 172 1998
rect 400 1964 448 1998
rect 676 1964 724 1998
rect 952 1964 1000 1998
rect 1228 1964 1276 1998
rect 1504 1964 1552 1998
rect 1780 1964 1828 1998
rect 2056 1964 2104 1998
rect 2332 1964 2380 1998
rect 2608 1964 2656 1998
rect 2884 1964 2932 1998
rect 3160 1964 3208 1998
rect 3436 1964 3484 1998
rect 3712 1964 3760 1998
rect 3988 1964 4036 1998
rect 4264 1964 4312 1998
rect 4540 1964 4588 1998
rect 4816 1964 4864 1998
rect 5092 1964 5140 1998
rect 5368 1964 5474 1998
rect 66 1952 5474 1964
rect 66 1902 124 1952
rect 66 1128 78 1902
rect 112 1128 124 1902
rect 5416 1902 5474 1952
rect 66 1078 124 1128
rect 5416 1128 5428 1902
rect 5462 1128 5474 1902
rect 5416 1078 5474 1128
rect 66 1066 5474 1078
rect 66 1032 172 1066
rect 400 1032 448 1066
rect 676 1032 724 1066
rect 952 1032 1000 1066
rect 1228 1032 1276 1066
rect 1504 1032 1552 1066
rect 1780 1032 1828 1066
rect 2056 1032 2104 1066
rect 2332 1032 2380 1066
rect 2608 1032 2656 1066
rect 2884 1032 2932 1066
rect 3160 1032 3208 1066
rect 3436 1032 3484 1066
rect 3712 1032 3760 1066
rect 3988 1032 4036 1066
rect 4264 1032 4312 1066
rect 4540 1032 4588 1066
rect 4816 1032 4864 1066
rect 5092 1032 5140 1066
rect 5368 1032 5474 1066
rect 66 1020 5474 1032
<< mvpsubdiffcont >>
rect 172 822 400 856
rect 448 822 676 856
rect 724 822 952 856
rect 1000 822 1228 856
rect 1276 822 1504 856
rect 1552 822 1780 856
rect 1828 822 2056 856
rect 2104 822 2332 856
rect 2380 822 2608 856
rect 2656 822 2884 856
rect 2932 822 3160 856
rect 3208 822 3436 856
rect 3484 822 3712 856
rect 3760 822 3988 856
rect 4036 822 4264 856
rect 4312 822 4540 856
rect 4588 822 4816 856
rect 4864 822 5092 856
rect 5140 822 5368 856
rect 58 144 92 760
rect 5458 144 5492 760
rect 172 48 400 82
rect 448 48 676 82
rect 724 48 952 82
rect 1000 48 1228 82
rect 1276 48 1504 82
rect 1552 48 1780 82
rect 1828 48 2056 82
rect 2104 48 2332 82
rect 2380 48 2608 82
rect 2656 48 2884 82
rect 2932 48 3160 82
rect 3208 48 3436 82
rect 3484 48 3712 82
rect 3760 48 3988 82
rect 4036 48 4264 82
rect 4312 48 4540 82
rect 4588 48 4816 82
rect 4864 48 5092 82
rect 5140 48 5368 82
<< mvnsubdiffcont >>
rect 172 1964 400 1998
rect 448 1964 676 1998
rect 724 1964 952 1998
rect 1000 1964 1228 1998
rect 1276 1964 1504 1998
rect 1552 1964 1780 1998
rect 1828 1964 2056 1998
rect 2104 1964 2332 1998
rect 2380 1964 2608 1998
rect 2656 1964 2884 1998
rect 2932 1964 3160 1998
rect 3208 1964 3436 1998
rect 3484 1964 3712 1998
rect 3760 1964 3988 1998
rect 4036 1964 4264 1998
rect 4312 1964 4540 1998
rect 4588 1964 4816 1998
rect 4864 1964 5092 1998
rect 5140 1964 5368 1998
rect 78 1128 112 1902
rect 5428 1128 5462 1902
rect 172 1032 400 1066
rect 448 1032 676 1066
rect 724 1032 952 1066
rect 1000 1032 1228 1066
rect 1276 1032 1504 1066
rect 1552 1032 1780 1066
rect 1828 1032 2056 1066
rect 2104 1032 2332 1066
rect 2380 1032 2608 1066
rect 2656 1032 2884 1066
rect 2932 1032 3160 1066
rect 3208 1032 3436 1066
rect 3484 1032 3712 1066
rect 3760 1032 3988 1066
rect 4036 1032 4264 1066
rect 4312 1032 4540 1066
rect 4588 1032 4816 1066
rect 4864 1032 5092 1066
rect 5140 1032 5368 1066
<< poly >>
rect 236 1914 336 1930
rect 236 1880 252 1914
rect 320 1880 336 1914
rect 236 1833 336 1880
rect 512 1914 612 1930
rect 512 1880 528 1914
rect 596 1880 612 1914
rect 512 1833 612 1880
rect 788 1914 888 1930
rect 788 1880 804 1914
rect 872 1880 888 1914
rect 788 1833 888 1880
rect 1064 1914 1164 1930
rect 1064 1880 1080 1914
rect 1148 1880 1164 1914
rect 1064 1833 1164 1880
rect 1340 1914 1440 1930
rect 1340 1880 1356 1914
rect 1424 1880 1440 1914
rect 1340 1833 1440 1880
rect 1616 1914 1716 1930
rect 1616 1880 1632 1914
rect 1700 1880 1716 1914
rect 1616 1833 1716 1880
rect 1892 1914 1992 1930
rect 1892 1880 1908 1914
rect 1976 1880 1992 1914
rect 1892 1833 1992 1880
rect 2168 1914 2268 1930
rect 2168 1880 2184 1914
rect 2252 1880 2268 1914
rect 2168 1833 2268 1880
rect 2444 1914 2544 1930
rect 2444 1880 2460 1914
rect 2528 1880 2544 1914
rect 2444 1833 2544 1880
rect 2720 1914 2820 1930
rect 2720 1880 2736 1914
rect 2804 1880 2820 1914
rect 2720 1833 2820 1880
rect 2996 1914 3096 1930
rect 2996 1880 3012 1914
rect 3080 1880 3096 1914
rect 2996 1833 3096 1880
rect 3272 1914 3372 1930
rect 3272 1880 3288 1914
rect 3356 1880 3372 1914
rect 3272 1833 3372 1880
rect 3548 1914 3648 1930
rect 3548 1880 3564 1914
rect 3632 1880 3648 1914
rect 3548 1833 3648 1880
rect 3824 1914 3924 1930
rect 3824 1880 3840 1914
rect 3908 1880 3924 1914
rect 3824 1833 3924 1880
rect 4100 1914 4200 1930
rect 4100 1880 4116 1914
rect 4184 1880 4200 1914
rect 4100 1833 4200 1880
rect 4376 1914 4476 1930
rect 4376 1880 4392 1914
rect 4460 1880 4476 1914
rect 4376 1833 4476 1880
rect 4652 1914 4752 1930
rect 4652 1880 4668 1914
rect 4736 1880 4752 1914
rect 4652 1833 4752 1880
rect 4928 1914 5028 1930
rect 4928 1880 4944 1914
rect 5012 1880 5028 1914
rect 4928 1833 5028 1880
rect 5204 1914 5304 1930
rect 5204 1880 5220 1914
rect 5288 1880 5304 1914
rect 5204 1833 5304 1880
rect 236 1586 336 1633
rect 236 1552 252 1586
rect 320 1552 336 1586
rect 236 1536 336 1552
rect 512 1586 612 1633
rect 512 1552 528 1586
rect 596 1552 612 1586
rect 512 1536 612 1552
rect 788 1586 888 1633
rect 788 1552 804 1586
rect 872 1552 888 1586
rect 788 1536 888 1552
rect 1064 1586 1164 1633
rect 1064 1552 1080 1586
rect 1148 1552 1164 1586
rect 1064 1536 1164 1552
rect 1340 1586 1440 1633
rect 1340 1552 1356 1586
rect 1424 1552 1440 1586
rect 1340 1536 1440 1552
rect 1616 1586 1716 1633
rect 1616 1552 1632 1586
rect 1700 1552 1716 1586
rect 1616 1536 1716 1552
rect 1892 1586 1992 1633
rect 1892 1552 1908 1586
rect 1976 1552 1992 1586
rect 1892 1536 1992 1552
rect 2168 1586 2268 1633
rect 2168 1552 2184 1586
rect 2252 1552 2268 1586
rect 2168 1536 2268 1552
rect 2444 1586 2544 1633
rect 2444 1552 2460 1586
rect 2528 1552 2544 1586
rect 2444 1536 2544 1552
rect 2720 1586 2820 1633
rect 2720 1552 2736 1586
rect 2804 1552 2820 1586
rect 2720 1536 2820 1552
rect 2996 1586 3096 1633
rect 2996 1552 3012 1586
rect 3080 1552 3096 1586
rect 2996 1536 3096 1552
rect 3272 1586 3372 1633
rect 3272 1552 3288 1586
rect 3356 1552 3372 1586
rect 3272 1536 3372 1552
rect 3548 1586 3648 1633
rect 3548 1552 3564 1586
rect 3632 1552 3648 1586
rect 3548 1536 3648 1552
rect 3824 1586 3924 1633
rect 3824 1552 3840 1586
rect 3908 1552 3924 1586
rect 3824 1536 3924 1552
rect 4100 1586 4200 1633
rect 4100 1552 4116 1586
rect 4184 1552 4200 1586
rect 4100 1536 4200 1552
rect 4376 1586 4476 1633
rect 4376 1552 4392 1586
rect 4460 1552 4476 1586
rect 4376 1536 4476 1552
rect 4652 1586 4752 1633
rect 4652 1552 4668 1586
rect 4736 1552 4752 1586
rect 4652 1536 4752 1552
rect 4928 1586 5028 1633
rect 4928 1552 4944 1586
rect 5012 1552 5028 1586
rect 4928 1536 5028 1552
rect 5204 1586 5304 1633
rect 5204 1552 5220 1586
rect 5288 1552 5304 1586
rect 5204 1536 5304 1552
rect 236 1478 336 1494
rect 236 1444 252 1478
rect 320 1444 336 1478
rect 236 1397 336 1444
rect 512 1478 612 1494
rect 512 1444 528 1478
rect 596 1444 612 1478
rect 512 1397 612 1444
rect 788 1478 888 1494
rect 788 1444 804 1478
rect 872 1444 888 1478
rect 788 1397 888 1444
rect 1064 1478 1164 1494
rect 1064 1444 1080 1478
rect 1148 1444 1164 1478
rect 1064 1397 1164 1444
rect 1340 1478 1440 1494
rect 1340 1444 1356 1478
rect 1424 1444 1440 1478
rect 1340 1397 1440 1444
rect 1616 1478 1716 1494
rect 1616 1444 1632 1478
rect 1700 1444 1716 1478
rect 1616 1397 1716 1444
rect 1892 1478 1992 1494
rect 1892 1444 1908 1478
rect 1976 1444 1992 1478
rect 1892 1397 1992 1444
rect 2168 1478 2268 1494
rect 2168 1444 2184 1478
rect 2252 1444 2268 1478
rect 2168 1397 2268 1444
rect 2444 1478 2544 1494
rect 2444 1444 2460 1478
rect 2528 1444 2544 1478
rect 2444 1397 2544 1444
rect 2720 1478 2820 1494
rect 2720 1444 2736 1478
rect 2804 1444 2820 1478
rect 2720 1397 2820 1444
rect 2996 1478 3096 1494
rect 2996 1444 3012 1478
rect 3080 1444 3096 1478
rect 2996 1397 3096 1444
rect 3272 1478 3372 1494
rect 3272 1444 3288 1478
rect 3356 1444 3372 1478
rect 3272 1397 3372 1444
rect 3548 1478 3648 1494
rect 3548 1444 3564 1478
rect 3632 1444 3648 1478
rect 3548 1397 3648 1444
rect 3824 1478 3924 1494
rect 3824 1444 3840 1478
rect 3908 1444 3924 1478
rect 3824 1397 3924 1444
rect 4100 1478 4200 1494
rect 4100 1444 4116 1478
rect 4184 1444 4200 1478
rect 4100 1397 4200 1444
rect 4376 1478 4476 1494
rect 4376 1444 4392 1478
rect 4460 1444 4476 1478
rect 4376 1397 4476 1444
rect 4652 1478 4752 1494
rect 4652 1444 4668 1478
rect 4736 1444 4752 1478
rect 4652 1397 4752 1444
rect 4928 1478 5028 1494
rect 4928 1444 4944 1478
rect 5012 1444 5028 1478
rect 4928 1397 5028 1444
rect 5204 1478 5304 1494
rect 5204 1444 5220 1478
rect 5288 1444 5304 1478
rect 5204 1397 5304 1444
rect 236 1150 336 1197
rect 236 1116 252 1150
rect 320 1116 336 1150
rect 236 1100 336 1116
rect 512 1150 612 1197
rect 512 1116 528 1150
rect 596 1116 612 1150
rect 512 1100 612 1116
rect 788 1150 888 1197
rect 788 1116 804 1150
rect 872 1116 888 1150
rect 788 1100 888 1116
rect 1064 1150 1164 1197
rect 1064 1116 1080 1150
rect 1148 1116 1164 1150
rect 1064 1100 1164 1116
rect 1340 1150 1440 1197
rect 1340 1116 1356 1150
rect 1424 1116 1440 1150
rect 1340 1100 1440 1116
rect 1616 1150 1716 1197
rect 1616 1116 1632 1150
rect 1700 1116 1716 1150
rect 1616 1100 1716 1116
rect 1892 1150 1992 1197
rect 1892 1116 1908 1150
rect 1976 1116 1992 1150
rect 1892 1100 1992 1116
rect 2168 1150 2268 1197
rect 2168 1116 2184 1150
rect 2252 1116 2268 1150
rect 2168 1100 2268 1116
rect 2444 1150 2544 1197
rect 2444 1116 2460 1150
rect 2528 1116 2544 1150
rect 2444 1100 2544 1116
rect 2720 1150 2820 1197
rect 2720 1116 2736 1150
rect 2804 1116 2820 1150
rect 2720 1100 2820 1116
rect 2996 1150 3096 1197
rect 2996 1116 3012 1150
rect 3080 1116 3096 1150
rect 2996 1100 3096 1116
rect 3272 1150 3372 1197
rect 3272 1116 3288 1150
rect 3356 1116 3372 1150
rect 3272 1100 3372 1116
rect 3548 1150 3648 1197
rect 3548 1116 3564 1150
rect 3632 1116 3648 1150
rect 3548 1100 3648 1116
rect 3824 1150 3924 1197
rect 3824 1116 3840 1150
rect 3908 1116 3924 1150
rect 3824 1100 3924 1116
rect 4100 1150 4200 1197
rect 4100 1116 4116 1150
rect 4184 1116 4200 1150
rect 4100 1100 4200 1116
rect 4376 1150 4476 1197
rect 4376 1116 4392 1150
rect 4460 1116 4476 1150
rect 4376 1100 4476 1116
rect 4652 1150 4752 1197
rect 4652 1116 4668 1150
rect 4736 1116 4752 1150
rect 4652 1100 4752 1116
rect 4928 1150 5028 1197
rect 4928 1116 4944 1150
rect 5012 1116 5028 1150
rect 4928 1100 5028 1116
rect 5204 1150 5304 1197
rect 5204 1116 5220 1150
rect 5288 1116 5304 1150
rect 5204 1100 5304 1116
rect 236 763 336 779
rect 236 729 252 763
rect 320 729 336 763
rect 236 691 336 729
rect 512 763 612 779
rect 512 729 528 763
rect 596 729 612 763
rect 512 691 612 729
rect 788 763 888 779
rect 788 729 804 763
rect 872 729 888 763
rect 788 691 888 729
rect 1064 763 1164 779
rect 1064 729 1080 763
rect 1148 729 1164 763
rect 1064 691 1164 729
rect 1340 763 1440 779
rect 1340 729 1356 763
rect 1424 729 1440 763
rect 1340 691 1440 729
rect 1616 763 1716 779
rect 1616 729 1632 763
rect 1700 729 1716 763
rect 1616 691 1716 729
rect 1892 763 1992 779
rect 1892 729 1908 763
rect 1976 729 1992 763
rect 1892 691 1992 729
rect 2168 763 2268 779
rect 2168 729 2184 763
rect 2252 729 2268 763
rect 2168 691 2268 729
rect 2444 763 2544 779
rect 2444 729 2460 763
rect 2528 729 2544 763
rect 2444 691 2544 729
rect 2720 763 2820 779
rect 2720 729 2736 763
rect 2804 729 2820 763
rect 2720 691 2820 729
rect 2996 763 3096 779
rect 2996 729 3012 763
rect 3080 729 3096 763
rect 2996 691 3096 729
rect 3272 763 3372 779
rect 3272 729 3288 763
rect 3356 729 3372 763
rect 3272 691 3372 729
rect 3548 763 3648 779
rect 3548 729 3564 763
rect 3632 729 3648 763
rect 3548 691 3648 729
rect 3824 763 3924 779
rect 3824 729 3840 763
rect 3908 729 3924 763
rect 3824 691 3924 729
rect 4100 763 4200 779
rect 4100 729 4116 763
rect 4184 729 4200 763
rect 4100 691 4200 729
rect 4376 763 4476 779
rect 4376 729 4392 763
rect 4460 729 4476 763
rect 4376 691 4476 729
rect 4652 763 4752 779
rect 4652 729 4668 763
rect 4736 729 4752 763
rect 4652 691 4752 729
rect 4928 763 5028 779
rect 4928 729 4944 763
rect 5012 729 5028 763
rect 4928 691 5028 729
rect 5204 763 5304 779
rect 5204 729 5220 763
rect 5288 729 5304 763
rect 5204 691 5304 729
rect 236 523 336 561
rect 236 489 252 523
rect 320 489 336 523
rect 236 473 336 489
rect 512 523 612 561
rect 512 489 528 523
rect 596 489 612 523
rect 512 473 612 489
rect 788 523 888 561
rect 788 489 804 523
rect 872 489 888 523
rect 788 473 888 489
rect 1064 523 1164 561
rect 1064 489 1080 523
rect 1148 489 1164 523
rect 1064 473 1164 489
rect 1340 523 1440 561
rect 1340 489 1356 523
rect 1424 489 1440 523
rect 1340 473 1440 489
rect 1616 523 1716 561
rect 1616 489 1632 523
rect 1700 489 1716 523
rect 1616 473 1716 489
rect 1892 523 1992 561
rect 1892 489 1908 523
rect 1976 489 1992 523
rect 1892 473 1992 489
rect 2168 523 2268 561
rect 2168 489 2184 523
rect 2252 489 2268 523
rect 2168 473 2268 489
rect 2444 523 2544 561
rect 2444 489 2460 523
rect 2528 489 2544 523
rect 2444 473 2544 489
rect 2720 523 2820 561
rect 2720 489 2736 523
rect 2804 489 2820 523
rect 2720 473 2820 489
rect 2996 523 3096 561
rect 2996 489 3012 523
rect 3080 489 3096 523
rect 2996 473 3096 489
rect 3272 523 3372 561
rect 3272 489 3288 523
rect 3356 489 3372 523
rect 3272 473 3372 489
rect 3548 523 3648 561
rect 3548 489 3564 523
rect 3632 489 3648 523
rect 3548 473 3648 489
rect 3824 523 3924 561
rect 3824 489 3840 523
rect 3908 489 3924 523
rect 3824 473 3924 489
rect 4100 523 4200 561
rect 4100 489 4116 523
rect 4184 489 4200 523
rect 4100 473 4200 489
rect 4376 523 4476 561
rect 4376 489 4392 523
rect 4460 489 4476 523
rect 4376 473 4476 489
rect 4652 523 4752 561
rect 4652 489 4668 523
rect 4736 489 4752 523
rect 4652 473 4752 489
rect 4928 523 5028 561
rect 4928 489 4944 523
rect 5012 489 5028 523
rect 4928 473 5028 489
rect 5204 523 5304 561
rect 5204 489 5220 523
rect 5288 489 5304 523
rect 5204 473 5304 489
rect 236 415 336 431
rect 236 381 252 415
rect 320 381 336 415
rect 236 343 336 381
rect 512 415 612 431
rect 512 381 528 415
rect 596 381 612 415
rect 512 343 612 381
rect 788 415 888 431
rect 788 381 804 415
rect 872 381 888 415
rect 788 343 888 381
rect 1064 415 1164 431
rect 1064 381 1080 415
rect 1148 381 1164 415
rect 1064 343 1164 381
rect 1340 415 1440 431
rect 1340 381 1356 415
rect 1424 381 1440 415
rect 1340 343 1440 381
rect 1616 415 1716 431
rect 1616 381 1632 415
rect 1700 381 1716 415
rect 1616 343 1716 381
rect 1892 415 1992 431
rect 1892 381 1908 415
rect 1976 381 1992 415
rect 1892 343 1992 381
rect 2168 415 2268 431
rect 2168 381 2184 415
rect 2252 381 2268 415
rect 2168 343 2268 381
rect 2444 415 2544 431
rect 2444 381 2460 415
rect 2528 381 2544 415
rect 2444 343 2544 381
rect 2720 415 2820 431
rect 2720 381 2736 415
rect 2804 381 2820 415
rect 2720 343 2820 381
rect 2996 415 3096 431
rect 2996 381 3012 415
rect 3080 381 3096 415
rect 2996 343 3096 381
rect 3272 415 3372 431
rect 3272 381 3288 415
rect 3356 381 3372 415
rect 3272 343 3372 381
rect 3548 415 3648 431
rect 3548 381 3564 415
rect 3632 381 3648 415
rect 3548 343 3648 381
rect 3824 415 3924 431
rect 3824 381 3840 415
rect 3908 381 3924 415
rect 3824 343 3924 381
rect 4100 415 4200 431
rect 4100 381 4116 415
rect 4184 381 4200 415
rect 4100 343 4200 381
rect 4376 415 4476 431
rect 4376 381 4392 415
rect 4460 381 4476 415
rect 4376 343 4476 381
rect 4652 415 4752 431
rect 4652 381 4668 415
rect 4736 381 4752 415
rect 4652 343 4752 381
rect 4928 415 5028 431
rect 4928 381 4944 415
rect 5012 381 5028 415
rect 4928 343 5028 381
rect 5204 415 5304 431
rect 5204 381 5220 415
rect 5288 381 5304 415
rect 5204 343 5304 381
rect 236 175 336 213
rect 236 141 252 175
rect 320 141 336 175
rect 236 125 336 141
rect 512 175 612 213
rect 512 141 528 175
rect 596 141 612 175
rect 512 125 612 141
rect 788 175 888 213
rect 788 141 804 175
rect 872 141 888 175
rect 788 125 888 141
rect 1064 175 1164 213
rect 1064 141 1080 175
rect 1148 141 1164 175
rect 1064 125 1164 141
rect 1340 175 1440 213
rect 1340 141 1356 175
rect 1424 141 1440 175
rect 1340 125 1440 141
rect 1616 175 1716 213
rect 1616 141 1632 175
rect 1700 141 1716 175
rect 1616 125 1716 141
rect 1892 175 1992 213
rect 1892 141 1908 175
rect 1976 141 1992 175
rect 1892 125 1992 141
rect 2168 175 2268 213
rect 2168 141 2184 175
rect 2252 141 2268 175
rect 2168 125 2268 141
rect 2444 175 2544 213
rect 2444 141 2460 175
rect 2528 141 2544 175
rect 2444 125 2544 141
rect 2720 175 2820 213
rect 2720 141 2736 175
rect 2804 141 2820 175
rect 2720 125 2820 141
rect 2996 175 3096 213
rect 2996 141 3012 175
rect 3080 141 3096 175
rect 2996 125 3096 141
rect 3272 175 3372 213
rect 3272 141 3288 175
rect 3356 141 3372 175
rect 3272 125 3372 141
rect 3548 175 3648 213
rect 3548 141 3564 175
rect 3632 141 3648 175
rect 3548 125 3648 141
rect 3824 175 3924 213
rect 3824 141 3840 175
rect 3908 141 3924 175
rect 3824 125 3924 141
rect 4100 175 4200 213
rect 4100 141 4116 175
rect 4184 141 4200 175
rect 4100 125 4200 141
rect 4376 175 4476 213
rect 4376 141 4392 175
rect 4460 141 4476 175
rect 4376 125 4476 141
rect 4652 175 4752 213
rect 4652 141 4668 175
rect 4736 141 4752 175
rect 4652 125 4752 141
rect 4928 175 5028 213
rect 4928 141 4944 175
rect 5012 141 5028 175
rect 4928 125 5028 141
rect 5204 175 5304 213
rect 5204 141 5220 175
rect 5288 141 5304 175
rect 5204 125 5304 141
<< polycont >>
rect 252 1880 320 1914
rect 528 1880 596 1914
rect 804 1880 872 1914
rect 1080 1880 1148 1914
rect 1356 1880 1424 1914
rect 1632 1880 1700 1914
rect 1908 1880 1976 1914
rect 2184 1880 2252 1914
rect 2460 1880 2528 1914
rect 2736 1880 2804 1914
rect 3012 1880 3080 1914
rect 3288 1880 3356 1914
rect 3564 1880 3632 1914
rect 3840 1880 3908 1914
rect 4116 1880 4184 1914
rect 4392 1880 4460 1914
rect 4668 1880 4736 1914
rect 4944 1880 5012 1914
rect 5220 1880 5288 1914
rect 252 1552 320 1586
rect 528 1552 596 1586
rect 804 1552 872 1586
rect 1080 1552 1148 1586
rect 1356 1552 1424 1586
rect 1632 1552 1700 1586
rect 1908 1552 1976 1586
rect 2184 1552 2252 1586
rect 2460 1552 2528 1586
rect 2736 1552 2804 1586
rect 3012 1552 3080 1586
rect 3288 1552 3356 1586
rect 3564 1552 3632 1586
rect 3840 1552 3908 1586
rect 4116 1552 4184 1586
rect 4392 1552 4460 1586
rect 4668 1552 4736 1586
rect 4944 1552 5012 1586
rect 5220 1552 5288 1586
rect 252 1444 320 1478
rect 528 1444 596 1478
rect 804 1444 872 1478
rect 1080 1444 1148 1478
rect 1356 1444 1424 1478
rect 1632 1444 1700 1478
rect 1908 1444 1976 1478
rect 2184 1444 2252 1478
rect 2460 1444 2528 1478
rect 2736 1444 2804 1478
rect 3012 1444 3080 1478
rect 3288 1444 3356 1478
rect 3564 1444 3632 1478
rect 3840 1444 3908 1478
rect 4116 1444 4184 1478
rect 4392 1444 4460 1478
rect 4668 1444 4736 1478
rect 4944 1444 5012 1478
rect 5220 1444 5288 1478
rect 252 1116 320 1150
rect 528 1116 596 1150
rect 804 1116 872 1150
rect 1080 1116 1148 1150
rect 1356 1116 1424 1150
rect 1632 1116 1700 1150
rect 1908 1116 1976 1150
rect 2184 1116 2252 1150
rect 2460 1116 2528 1150
rect 2736 1116 2804 1150
rect 3012 1116 3080 1150
rect 3288 1116 3356 1150
rect 3564 1116 3632 1150
rect 3840 1116 3908 1150
rect 4116 1116 4184 1150
rect 4392 1116 4460 1150
rect 4668 1116 4736 1150
rect 4944 1116 5012 1150
rect 5220 1116 5288 1150
rect 252 729 320 763
rect 528 729 596 763
rect 804 729 872 763
rect 1080 729 1148 763
rect 1356 729 1424 763
rect 1632 729 1700 763
rect 1908 729 1976 763
rect 2184 729 2252 763
rect 2460 729 2528 763
rect 2736 729 2804 763
rect 3012 729 3080 763
rect 3288 729 3356 763
rect 3564 729 3632 763
rect 3840 729 3908 763
rect 4116 729 4184 763
rect 4392 729 4460 763
rect 4668 729 4736 763
rect 4944 729 5012 763
rect 5220 729 5288 763
rect 252 489 320 523
rect 528 489 596 523
rect 804 489 872 523
rect 1080 489 1148 523
rect 1356 489 1424 523
rect 1632 489 1700 523
rect 1908 489 1976 523
rect 2184 489 2252 523
rect 2460 489 2528 523
rect 2736 489 2804 523
rect 3012 489 3080 523
rect 3288 489 3356 523
rect 3564 489 3632 523
rect 3840 489 3908 523
rect 4116 489 4184 523
rect 4392 489 4460 523
rect 4668 489 4736 523
rect 4944 489 5012 523
rect 5220 489 5288 523
rect 252 381 320 415
rect 528 381 596 415
rect 804 381 872 415
rect 1080 381 1148 415
rect 1356 381 1424 415
rect 1632 381 1700 415
rect 1908 381 1976 415
rect 2184 381 2252 415
rect 2460 381 2528 415
rect 2736 381 2804 415
rect 3012 381 3080 415
rect 3288 381 3356 415
rect 3564 381 3632 415
rect 3840 381 3908 415
rect 4116 381 4184 415
rect 4392 381 4460 415
rect 4668 381 4736 415
rect 4944 381 5012 415
rect 5220 381 5288 415
rect 252 141 320 175
rect 528 141 596 175
rect 804 141 872 175
rect 1080 141 1148 175
rect 1356 141 1424 175
rect 1632 141 1700 175
rect 1908 141 1976 175
rect 2184 141 2252 175
rect 2460 141 2528 175
rect 2736 141 2804 175
rect 3012 141 3080 175
rect 3288 141 3356 175
rect 3564 141 3632 175
rect 3840 141 3908 175
rect 4116 141 4184 175
rect 4392 141 4460 175
rect 4668 141 4736 175
rect 4944 141 5012 175
rect 5220 141 5288 175
<< locali >>
rect 78 1964 172 1998
rect 400 1964 448 1998
rect 676 1964 724 1998
rect 952 1964 1000 1998
rect 1228 1964 1276 1998
rect 1504 1964 1552 1998
rect 1780 1964 1828 1998
rect 2056 1964 2104 1998
rect 2332 1964 2380 1998
rect 2608 1964 2656 1998
rect 2884 1964 2932 1998
rect 3160 1964 3208 1998
rect 3436 1964 3484 1998
rect 3712 1964 3760 1998
rect 3988 1964 4036 1998
rect 4264 1964 4312 1998
rect 4540 1964 4588 1998
rect 4816 1964 4864 1998
rect 5092 1964 5140 1998
rect 5368 1964 5462 1998
rect 78 1902 112 1964
rect 236 1880 252 1914
rect 320 1880 336 1914
rect 512 1880 528 1914
rect 596 1880 612 1914
rect 788 1880 804 1914
rect 872 1880 888 1914
rect 1064 1880 1080 1914
rect 1148 1880 1164 1914
rect 1340 1880 1356 1914
rect 1424 1880 1440 1914
rect 1616 1880 1632 1914
rect 1700 1880 1716 1914
rect 1892 1880 1908 1914
rect 1976 1880 1992 1914
rect 2168 1880 2184 1914
rect 2252 1880 2268 1914
rect 2444 1880 2460 1914
rect 2528 1880 2544 1914
rect 2720 1880 2736 1914
rect 2804 1880 2820 1914
rect 2996 1880 3012 1914
rect 3080 1880 3096 1914
rect 3272 1880 3288 1914
rect 3356 1880 3372 1914
rect 3548 1880 3564 1914
rect 3632 1880 3648 1914
rect 3824 1880 3840 1914
rect 3908 1880 3924 1914
rect 4100 1880 4116 1914
rect 4184 1880 4200 1914
rect 4376 1880 4392 1914
rect 4460 1880 4476 1914
rect 4652 1880 4668 1914
rect 4736 1880 4752 1914
rect 4928 1880 4944 1914
rect 5012 1880 5028 1914
rect 5204 1880 5220 1914
rect 5288 1880 5304 1914
rect 5428 1902 5462 1964
rect 190 1821 224 1837
rect 190 1629 224 1645
rect 348 1821 382 1837
rect 348 1629 382 1645
rect 466 1821 500 1837
rect 466 1629 500 1645
rect 624 1821 658 1837
rect 624 1629 658 1645
rect 742 1821 776 1837
rect 742 1629 776 1645
rect 900 1821 934 1837
rect 900 1629 934 1645
rect 1018 1821 1052 1837
rect 1018 1629 1052 1645
rect 1176 1821 1210 1837
rect 1176 1629 1210 1645
rect 1294 1821 1328 1837
rect 1294 1629 1328 1645
rect 1452 1821 1486 1837
rect 1452 1629 1486 1645
rect 1570 1821 1604 1837
rect 1570 1629 1604 1645
rect 1728 1821 1762 1837
rect 1728 1629 1762 1645
rect 1846 1821 1880 1837
rect 1846 1629 1880 1645
rect 2004 1821 2038 1837
rect 2004 1629 2038 1645
rect 2122 1821 2156 1837
rect 2122 1629 2156 1645
rect 2280 1821 2314 1837
rect 2280 1629 2314 1645
rect 2398 1821 2432 1837
rect 2398 1629 2432 1645
rect 2556 1821 2590 1837
rect 2556 1629 2590 1645
rect 2674 1821 2708 1837
rect 2674 1629 2708 1645
rect 2832 1821 2866 1837
rect 2832 1629 2866 1645
rect 2950 1821 2984 1837
rect 2950 1629 2984 1645
rect 3108 1821 3142 1837
rect 3108 1629 3142 1645
rect 3226 1821 3260 1837
rect 3226 1629 3260 1645
rect 3384 1821 3418 1837
rect 3384 1629 3418 1645
rect 3502 1821 3536 1837
rect 3502 1629 3536 1645
rect 3660 1821 3694 1837
rect 3660 1629 3694 1645
rect 3778 1821 3812 1837
rect 3778 1629 3812 1645
rect 3936 1821 3970 1837
rect 3936 1629 3970 1645
rect 4054 1821 4088 1837
rect 4054 1629 4088 1645
rect 4212 1821 4246 1837
rect 4212 1629 4246 1645
rect 4330 1821 4364 1837
rect 4330 1629 4364 1645
rect 4488 1821 4522 1837
rect 4488 1629 4522 1645
rect 4606 1821 4640 1837
rect 4606 1629 4640 1645
rect 4764 1821 4798 1837
rect 4764 1629 4798 1645
rect 4882 1821 4916 1837
rect 4882 1629 4916 1645
rect 5040 1821 5074 1837
rect 5040 1629 5074 1645
rect 5158 1821 5192 1837
rect 5158 1629 5192 1645
rect 5316 1821 5350 1837
rect 5316 1629 5350 1645
rect 236 1552 252 1586
rect 320 1552 336 1586
rect 512 1552 528 1586
rect 596 1552 612 1586
rect 788 1552 804 1586
rect 872 1552 888 1586
rect 1064 1552 1080 1586
rect 1148 1552 1164 1586
rect 1340 1552 1356 1586
rect 1424 1552 1440 1586
rect 1616 1552 1632 1586
rect 1700 1552 1716 1586
rect 1892 1552 1908 1586
rect 1976 1552 1992 1586
rect 2168 1552 2184 1586
rect 2252 1552 2268 1586
rect 2444 1552 2460 1586
rect 2528 1552 2544 1586
rect 2720 1552 2736 1586
rect 2804 1552 2820 1586
rect 2996 1552 3012 1586
rect 3080 1552 3096 1586
rect 3272 1552 3288 1586
rect 3356 1552 3372 1586
rect 3548 1552 3564 1586
rect 3632 1552 3648 1586
rect 3824 1552 3840 1586
rect 3908 1552 3924 1586
rect 4100 1552 4116 1586
rect 4184 1552 4200 1586
rect 4376 1552 4392 1586
rect 4460 1552 4476 1586
rect 4652 1552 4668 1586
rect 4736 1552 4752 1586
rect 4928 1552 4944 1586
rect 5012 1552 5028 1586
rect 5204 1552 5220 1586
rect 5288 1552 5304 1586
rect 236 1444 252 1478
rect 320 1444 336 1478
rect 512 1444 528 1478
rect 596 1444 612 1478
rect 788 1444 804 1478
rect 872 1444 888 1478
rect 1064 1444 1080 1478
rect 1148 1444 1164 1478
rect 1340 1444 1356 1478
rect 1424 1444 1440 1478
rect 1616 1444 1632 1478
rect 1700 1444 1716 1478
rect 1892 1444 1908 1478
rect 1976 1444 1992 1478
rect 2168 1444 2184 1478
rect 2252 1444 2268 1478
rect 2444 1444 2460 1478
rect 2528 1444 2544 1478
rect 2720 1444 2736 1478
rect 2804 1444 2820 1478
rect 2996 1444 3012 1478
rect 3080 1444 3096 1478
rect 3272 1444 3288 1478
rect 3356 1444 3372 1478
rect 3548 1444 3564 1478
rect 3632 1444 3648 1478
rect 3824 1444 3840 1478
rect 3908 1444 3924 1478
rect 4100 1444 4116 1478
rect 4184 1444 4200 1478
rect 4376 1444 4392 1478
rect 4460 1444 4476 1478
rect 4652 1444 4668 1478
rect 4736 1444 4752 1478
rect 4928 1444 4944 1478
rect 5012 1444 5028 1478
rect 5204 1444 5220 1478
rect 5288 1444 5304 1478
rect 190 1385 224 1401
rect 190 1193 224 1209
rect 348 1385 382 1401
rect 348 1193 382 1209
rect 466 1385 500 1401
rect 466 1193 500 1209
rect 624 1385 658 1401
rect 624 1193 658 1209
rect 742 1385 776 1401
rect 742 1193 776 1209
rect 900 1385 934 1401
rect 900 1193 934 1209
rect 1018 1385 1052 1401
rect 1018 1193 1052 1209
rect 1176 1385 1210 1401
rect 1176 1193 1210 1209
rect 1294 1385 1328 1401
rect 1294 1193 1328 1209
rect 1452 1385 1486 1401
rect 1452 1193 1486 1209
rect 1570 1385 1604 1401
rect 1570 1193 1604 1209
rect 1728 1385 1762 1401
rect 1728 1193 1762 1209
rect 1846 1385 1880 1401
rect 1846 1193 1880 1209
rect 2004 1385 2038 1401
rect 2004 1193 2038 1209
rect 2122 1385 2156 1401
rect 2122 1193 2156 1209
rect 2280 1385 2314 1401
rect 2280 1193 2314 1209
rect 2398 1385 2432 1401
rect 2398 1193 2432 1209
rect 2556 1385 2590 1401
rect 2556 1193 2590 1209
rect 2674 1385 2708 1401
rect 2674 1193 2708 1209
rect 2832 1385 2866 1401
rect 2832 1193 2866 1209
rect 2950 1385 2984 1401
rect 2950 1193 2984 1209
rect 3108 1385 3142 1401
rect 3108 1193 3142 1209
rect 3226 1385 3260 1401
rect 3226 1193 3260 1209
rect 3384 1385 3418 1401
rect 3384 1193 3418 1209
rect 3502 1385 3536 1401
rect 3502 1193 3536 1209
rect 3660 1385 3694 1401
rect 3660 1193 3694 1209
rect 3778 1385 3812 1401
rect 3778 1193 3812 1209
rect 3936 1385 3970 1401
rect 3936 1193 3970 1209
rect 4054 1385 4088 1401
rect 4054 1193 4088 1209
rect 4212 1385 4246 1401
rect 4212 1193 4246 1209
rect 4330 1385 4364 1401
rect 4330 1193 4364 1209
rect 4488 1385 4522 1401
rect 4488 1193 4522 1209
rect 4606 1385 4640 1401
rect 4606 1193 4640 1209
rect 4764 1385 4798 1401
rect 4764 1193 4798 1209
rect 4882 1385 4916 1401
rect 4882 1193 4916 1209
rect 5040 1385 5074 1401
rect 5040 1193 5074 1209
rect 5158 1385 5192 1401
rect 5158 1193 5192 1209
rect 5316 1385 5350 1401
rect 5316 1193 5350 1209
rect 78 1066 112 1128
rect 236 1116 252 1150
rect 320 1116 336 1150
rect 512 1116 528 1150
rect 596 1116 612 1150
rect 788 1116 804 1150
rect 872 1116 888 1150
rect 1064 1116 1080 1150
rect 1148 1116 1164 1150
rect 1340 1116 1356 1150
rect 1424 1116 1440 1150
rect 1616 1116 1632 1150
rect 1700 1116 1716 1150
rect 1892 1116 1908 1150
rect 1976 1116 1992 1150
rect 2168 1116 2184 1150
rect 2252 1116 2268 1150
rect 2444 1116 2460 1150
rect 2528 1116 2544 1150
rect 2720 1116 2736 1150
rect 2804 1116 2820 1150
rect 2996 1116 3012 1150
rect 3080 1116 3096 1150
rect 3272 1116 3288 1150
rect 3356 1116 3372 1150
rect 3548 1116 3564 1150
rect 3632 1116 3648 1150
rect 3824 1116 3840 1150
rect 3908 1116 3924 1150
rect 4100 1116 4116 1150
rect 4184 1116 4200 1150
rect 4376 1116 4392 1150
rect 4460 1116 4476 1150
rect 4652 1116 4668 1150
rect 4736 1116 4752 1150
rect 4928 1116 4944 1150
rect 5012 1116 5028 1150
rect 5204 1116 5220 1150
rect 5288 1116 5304 1150
rect 5428 1066 5462 1128
rect 78 1032 172 1066
rect 400 1032 448 1066
rect 676 1032 724 1066
rect 952 1032 1000 1066
rect 1228 1032 1276 1066
rect 1504 1032 1552 1066
rect 1780 1032 1828 1066
rect 2056 1032 2104 1066
rect 2332 1032 2380 1066
rect 2608 1032 2656 1066
rect 2884 1032 2932 1066
rect 3160 1032 3208 1066
rect 3436 1032 3484 1066
rect 3712 1032 3760 1066
rect 3988 1032 4036 1066
rect 4264 1032 4312 1066
rect 4540 1032 4588 1066
rect 4816 1032 4864 1066
rect 5092 1032 5140 1066
rect 5368 1032 5462 1066
rect 58 822 172 856
rect 400 822 448 856
rect 676 822 724 856
rect 952 822 1000 856
rect 1228 822 1276 856
rect 1504 822 1552 856
rect 1780 822 1828 856
rect 2056 822 2104 856
rect 2332 822 2380 856
rect 2608 822 2656 856
rect 2884 822 2932 856
rect 3160 822 3208 856
rect 3436 822 3484 856
rect 3712 822 3760 856
rect 3988 822 4036 856
rect 4264 822 4312 856
rect 4540 822 4588 856
rect 4816 822 4864 856
rect 5092 822 5140 856
rect 5368 822 5492 856
rect 58 760 92 822
rect 236 729 252 763
rect 320 729 336 763
rect 512 729 528 763
rect 596 729 612 763
rect 788 729 804 763
rect 872 729 888 763
rect 1064 729 1080 763
rect 1148 729 1164 763
rect 1340 729 1356 763
rect 1424 729 1440 763
rect 1616 729 1632 763
rect 1700 729 1716 763
rect 1892 729 1908 763
rect 1976 729 1992 763
rect 2168 729 2184 763
rect 2252 729 2268 763
rect 2444 729 2460 763
rect 2528 729 2544 763
rect 2720 729 2736 763
rect 2804 729 2820 763
rect 2996 729 3012 763
rect 3080 729 3096 763
rect 3272 729 3288 763
rect 3356 729 3372 763
rect 3548 729 3564 763
rect 3632 729 3648 763
rect 3824 729 3840 763
rect 3908 729 3924 763
rect 4100 729 4116 763
rect 4184 729 4200 763
rect 4376 729 4392 763
rect 4460 729 4476 763
rect 4652 729 4668 763
rect 4736 729 4752 763
rect 4928 729 4944 763
rect 5012 729 5028 763
rect 5204 729 5220 763
rect 5288 729 5304 763
rect 5458 760 5492 822
rect 190 679 224 695
rect 190 557 224 573
rect 348 679 382 695
rect 348 557 382 573
rect 466 679 500 695
rect 466 557 500 573
rect 624 679 658 695
rect 624 557 658 573
rect 742 679 776 695
rect 742 557 776 573
rect 900 679 934 695
rect 900 557 934 573
rect 1018 679 1052 695
rect 1018 557 1052 573
rect 1176 679 1210 695
rect 1176 557 1210 573
rect 1294 679 1328 695
rect 1294 557 1328 573
rect 1452 679 1486 695
rect 1452 557 1486 573
rect 1570 679 1604 695
rect 1570 557 1604 573
rect 1728 679 1762 695
rect 1728 557 1762 573
rect 1846 679 1880 695
rect 1846 557 1880 573
rect 2004 679 2038 695
rect 2004 557 2038 573
rect 2122 679 2156 695
rect 2122 557 2156 573
rect 2280 679 2314 695
rect 2280 557 2314 573
rect 2398 679 2432 695
rect 2398 557 2432 573
rect 2556 679 2590 695
rect 2556 557 2590 573
rect 2674 679 2708 695
rect 2674 557 2708 573
rect 2832 679 2866 695
rect 2832 557 2866 573
rect 2950 679 2984 695
rect 2950 557 2984 573
rect 3108 679 3142 695
rect 3108 557 3142 573
rect 3226 679 3260 695
rect 3226 557 3260 573
rect 3384 679 3418 695
rect 3384 557 3418 573
rect 3502 679 3536 695
rect 3502 557 3536 573
rect 3660 679 3694 695
rect 3660 557 3694 573
rect 3778 679 3812 695
rect 3778 557 3812 573
rect 3936 679 3970 695
rect 3936 557 3970 573
rect 4054 679 4088 695
rect 4054 557 4088 573
rect 4212 679 4246 695
rect 4212 557 4246 573
rect 4330 679 4364 695
rect 4330 557 4364 573
rect 4488 679 4522 695
rect 4488 557 4522 573
rect 4606 679 4640 695
rect 4606 557 4640 573
rect 4764 679 4798 695
rect 4764 557 4798 573
rect 4882 679 4916 695
rect 4882 557 4916 573
rect 5040 679 5074 695
rect 5040 557 5074 573
rect 5158 679 5192 695
rect 5158 557 5192 573
rect 5316 679 5350 695
rect 5316 557 5350 573
rect 236 489 252 523
rect 320 489 336 523
rect 512 489 528 523
rect 596 489 612 523
rect 788 489 804 523
rect 872 489 888 523
rect 1064 489 1080 523
rect 1148 489 1164 523
rect 1340 489 1356 523
rect 1424 489 1440 523
rect 1616 489 1632 523
rect 1700 489 1716 523
rect 1892 489 1908 523
rect 1976 489 1992 523
rect 2168 489 2184 523
rect 2252 489 2268 523
rect 2444 489 2460 523
rect 2528 489 2544 523
rect 2720 489 2736 523
rect 2804 489 2820 523
rect 2996 489 3012 523
rect 3080 489 3096 523
rect 3272 489 3288 523
rect 3356 489 3372 523
rect 3548 489 3564 523
rect 3632 489 3648 523
rect 3824 489 3840 523
rect 3908 489 3924 523
rect 4100 489 4116 523
rect 4184 489 4200 523
rect 4376 489 4392 523
rect 4460 489 4476 523
rect 4652 489 4668 523
rect 4736 489 4752 523
rect 4928 489 4944 523
rect 5012 489 5028 523
rect 5204 489 5220 523
rect 5288 489 5304 523
rect 236 381 252 415
rect 320 381 336 415
rect 512 381 528 415
rect 596 381 612 415
rect 788 381 804 415
rect 872 381 888 415
rect 1064 381 1080 415
rect 1148 381 1164 415
rect 1340 381 1356 415
rect 1424 381 1440 415
rect 1616 381 1632 415
rect 1700 381 1716 415
rect 1892 381 1908 415
rect 1976 381 1992 415
rect 2168 381 2184 415
rect 2252 381 2268 415
rect 2444 381 2460 415
rect 2528 381 2544 415
rect 2720 381 2736 415
rect 2804 381 2820 415
rect 2996 381 3012 415
rect 3080 381 3096 415
rect 3272 381 3288 415
rect 3356 381 3372 415
rect 3548 381 3564 415
rect 3632 381 3648 415
rect 3824 381 3840 415
rect 3908 381 3924 415
rect 4100 381 4116 415
rect 4184 381 4200 415
rect 4376 381 4392 415
rect 4460 381 4476 415
rect 4652 381 4668 415
rect 4736 381 4752 415
rect 4928 381 4944 415
rect 5012 381 5028 415
rect 5204 381 5220 415
rect 5288 381 5304 415
rect 190 331 224 347
rect 190 209 224 225
rect 348 331 382 347
rect 348 209 382 225
rect 466 331 500 347
rect 466 209 500 225
rect 624 331 658 347
rect 624 209 658 225
rect 742 331 776 347
rect 742 209 776 225
rect 900 331 934 347
rect 900 209 934 225
rect 1018 331 1052 347
rect 1018 209 1052 225
rect 1176 331 1210 347
rect 1176 209 1210 225
rect 1294 331 1328 347
rect 1294 209 1328 225
rect 1452 331 1486 347
rect 1452 209 1486 225
rect 1570 331 1604 347
rect 1570 209 1604 225
rect 1728 331 1762 347
rect 1728 209 1762 225
rect 1846 331 1880 347
rect 1846 209 1880 225
rect 2004 331 2038 347
rect 2004 209 2038 225
rect 2122 331 2156 347
rect 2122 209 2156 225
rect 2280 331 2314 347
rect 2280 209 2314 225
rect 2398 331 2432 347
rect 2398 209 2432 225
rect 2556 331 2590 347
rect 2556 209 2590 225
rect 2674 331 2708 347
rect 2674 209 2708 225
rect 2832 331 2866 347
rect 2832 209 2866 225
rect 2950 331 2984 347
rect 2950 209 2984 225
rect 3108 331 3142 347
rect 3108 209 3142 225
rect 3226 331 3260 347
rect 3226 209 3260 225
rect 3384 331 3418 347
rect 3384 209 3418 225
rect 3502 331 3536 347
rect 3502 209 3536 225
rect 3660 331 3694 347
rect 3660 209 3694 225
rect 3778 331 3812 347
rect 3778 209 3812 225
rect 3936 331 3970 347
rect 3936 209 3970 225
rect 4054 331 4088 347
rect 4054 209 4088 225
rect 4212 331 4246 347
rect 4212 209 4246 225
rect 4330 331 4364 347
rect 4330 209 4364 225
rect 4488 331 4522 347
rect 4488 209 4522 225
rect 4606 331 4640 347
rect 4606 209 4640 225
rect 4764 331 4798 347
rect 4764 209 4798 225
rect 4882 331 4916 347
rect 4882 209 4916 225
rect 5040 331 5074 347
rect 5040 209 5074 225
rect 5158 331 5192 347
rect 5158 209 5192 225
rect 5316 331 5350 347
rect 5316 209 5350 225
rect 58 82 92 144
rect 236 141 252 175
rect 320 141 336 175
rect 512 141 528 175
rect 596 141 612 175
rect 788 141 804 175
rect 872 141 888 175
rect 1064 141 1080 175
rect 1148 141 1164 175
rect 1340 141 1356 175
rect 1424 141 1440 175
rect 1616 141 1632 175
rect 1700 141 1716 175
rect 1892 141 1908 175
rect 1976 141 1992 175
rect 2168 141 2184 175
rect 2252 141 2268 175
rect 2444 141 2460 175
rect 2528 141 2544 175
rect 2720 141 2736 175
rect 2804 141 2820 175
rect 2996 141 3012 175
rect 3080 141 3096 175
rect 3272 141 3288 175
rect 3356 141 3372 175
rect 3548 141 3564 175
rect 3632 141 3648 175
rect 3824 141 3840 175
rect 3908 141 3924 175
rect 4100 141 4116 175
rect 4184 141 4200 175
rect 4376 141 4392 175
rect 4460 141 4476 175
rect 4652 141 4668 175
rect 4736 141 4752 175
rect 4928 141 4944 175
rect 5012 141 5028 175
rect 5204 141 5220 175
rect 5288 141 5304 175
rect 5458 82 5492 144
rect 58 48 172 82
rect 400 48 448 82
rect 676 48 724 82
rect 952 48 1000 82
rect 1228 48 1276 82
rect 1504 48 1552 82
rect 1780 48 1828 82
rect 2056 48 2104 82
rect 2332 48 2380 82
rect 2608 48 2656 82
rect 2884 48 2932 82
rect 3160 48 3208 82
rect 3436 48 3484 82
rect 3712 48 3760 82
rect 3988 48 4036 82
rect 4264 48 4312 82
rect 4540 48 4588 82
rect 4816 48 4864 82
rect 5092 48 5140 82
rect 5368 48 5492 82
<< viali >>
rect 172 1964 400 1998
rect 448 1964 676 1998
rect 724 1964 952 1998
rect 1000 1964 1228 1998
rect 1276 1964 1504 1998
rect 1552 1964 1780 1998
rect 1828 1964 2056 1998
rect 2104 1964 2332 1998
rect 2380 1964 2608 1998
rect 2656 1964 2884 1998
rect 2932 1964 3160 1998
rect 3208 1964 3436 1998
rect 3484 1964 3712 1998
rect 3760 1964 3988 1998
rect 4036 1964 4264 1998
rect 4312 1964 4540 1998
rect 4588 1964 4816 1998
rect 4864 1964 5092 1998
rect 5140 1964 5368 1998
rect 252 1880 320 1914
rect 528 1880 596 1914
rect 804 1880 872 1914
rect 1080 1880 1148 1914
rect 1356 1880 1424 1914
rect 1632 1880 1700 1914
rect 1908 1880 1976 1914
rect 2184 1880 2252 1914
rect 2460 1880 2528 1914
rect 2736 1880 2804 1914
rect 3012 1880 3080 1914
rect 3288 1880 3356 1914
rect 3564 1880 3632 1914
rect 3840 1880 3908 1914
rect 4116 1880 4184 1914
rect 4392 1880 4460 1914
rect 4668 1880 4736 1914
rect 4944 1880 5012 1914
rect 5220 1880 5288 1914
rect 190 1645 224 1821
rect 348 1645 382 1821
rect 466 1645 500 1821
rect 624 1645 658 1821
rect 742 1645 776 1821
rect 900 1645 934 1821
rect 1018 1645 1052 1821
rect 1176 1645 1210 1821
rect 1294 1645 1328 1821
rect 1452 1645 1486 1821
rect 1570 1645 1604 1821
rect 1728 1645 1762 1821
rect 1846 1645 1880 1821
rect 2004 1645 2038 1821
rect 2122 1645 2156 1821
rect 2280 1645 2314 1821
rect 2398 1645 2432 1821
rect 2556 1645 2590 1821
rect 2674 1645 2708 1821
rect 2832 1645 2866 1821
rect 2950 1645 2984 1821
rect 3108 1645 3142 1821
rect 3226 1645 3260 1821
rect 3384 1645 3418 1821
rect 3502 1645 3536 1821
rect 3660 1645 3694 1821
rect 3778 1645 3812 1821
rect 3936 1645 3970 1821
rect 4054 1645 4088 1821
rect 4212 1645 4246 1821
rect 4330 1645 4364 1821
rect 4488 1645 4522 1821
rect 4606 1645 4640 1821
rect 4764 1645 4798 1821
rect 4882 1645 4916 1821
rect 5040 1645 5074 1821
rect 5158 1645 5192 1821
rect 5316 1645 5350 1821
rect 252 1552 320 1586
rect 528 1552 596 1586
rect 804 1552 872 1586
rect 1080 1552 1148 1586
rect 1356 1552 1424 1586
rect 1632 1552 1700 1586
rect 1908 1552 1976 1586
rect 2184 1552 2252 1586
rect 2460 1552 2528 1586
rect 2736 1552 2804 1586
rect 3012 1552 3080 1586
rect 3288 1552 3356 1586
rect 3564 1552 3632 1586
rect 3840 1552 3908 1586
rect 4116 1552 4184 1586
rect 4392 1552 4460 1586
rect 4668 1552 4736 1586
rect 4944 1552 5012 1586
rect 5220 1552 5288 1586
rect 252 1444 320 1478
rect 528 1444 596 1478
rect 804 1444 872 1478
rect 1080 1444 1148 1478
rect 1356 1444 1424 1478
rect 1632 1444 1700 1478
rect 1908 1444 1976 1478
rect 2184 1444 2252 1478
rect 2460 1444 2528 1478
rect 2736 1444 2804 1478
rect 3012 1444 3080 1478
rect 3288 1444 3356 1478
rect 3564 1444 3632 1478
rect 3840 1444 3908 1478
rect 4116 1444 4184 1478
rect 4392 1444 4460 1478
rect 4668 1444 4736 1478
rect 4944 1444 5012 1478
rect 5220 1444 5288 1478
rect 190 1209 224 1385
rect 348 1209 382 1385
rect 466 1209 500 1385
rect 624 1209 658 1385
rect 742 1209 776 1385
rect 900 1209 934 1385
rect 1018 1209 1052 1385
rect 1176 1209 1210 1385
rect 1294 1209 1328 1385
rect 1452 1209 1486 1385
rect 1570 1209 1604 1385
rect 1728 1209 1762 1385
rect 1846 1209 1880 1385
rect 2004 1209 2038 1385
rect 2122 1209 2156 1385
rect 2280 1209 2314 1385
rect 2398 1209 2432 1385
rect 2556 1209 2590 1385
rect 2674 1209 2708 1385
rect 2832 1209 2866 1385
rect 2950 1209 2984 1385
rect 3108 1209 3142 1385
rect 3226 1209 3260 1385
rect 3384 1209 3418 1385
rect 3502 1209 3536 1385
rect 3660 1209 3694 1385
rect 3778 1209 3812 1385
rect 3936 1209 3970 1385
rect 4054 1209 4088 1385
rect 4212 1209 4246 1385
rect 4330 1209 4364 1385
rect 4488 1209 4522 1385
rect 4606 1209 4640 1385
rect 4764 1209 4798 1385
rect 4882 1209 4916 1385
rect 5040 1209 5074 1385
rect 5158 1209 5192 1385
rect 5316 1209 5350 1385
rect 252 1116 320 1150
rect 528 1116 596 1150
rect 804 1116 872 1150
rect 1080 1116 1148 1150
rect 1356 1116 1424 1150
rect 1632 1116 1700 1150
rect 1908 1116 1976 1150
rect 2184 1116 2252 1150
rect 2460 1116 2528 1150
rect 2736 1116 2804 1150
rect 3012 1116 3080 1150
rect 3288 1116 3356 1150
rect 3564 1116 3632 1150
rect 3840 1116 3908 1150
rect 4116 1116 4184 1150
rect 4392 1116 4460 1150
rect 4668 1116 4736 1150
rect 4944 1116 5012 1150
rect 5220 1116 5288 1150
rect 252 729 320 763
rect 528 729 596 763
rect 804 729 872 763
rect 1080 729 1148 763
rect 1356 729 1424 763
rect 1632 729 1700 763
rect 1908 729 1976 763
rect 2184 729 2252 763
rect 2460 729 2528 763
rect 2736 729 2804 763
rect 3012 729 3080 763
rect 3288 729 3356 763
rect 3564 729 3632 763
rect 3840 729 3908 763
rect 4116 729 4184 763
rect 4392 729 4460 763
rect 4668 729 4736 763
rect 4944 729 5012 763
rect 5220 729 5288 763
rect 190 573 224 679
rect 348 573 382 679
rect 466 573 500 679
rect 624 573 658 679
rect 742 573 776 679
rect 900 573 934 679
rect 1018 573 1052 679
rect 1176 573 1210 679
rect 1294 573 1328 679
rect 1452 573 1486 679
rect 1570 573 1604 679
rect 1728 573 1762 679
rect 1846 573 1880 679
rect 2004 573 2038 679
rect 2122 573 2156 679
rect 2280 573 2314 679
rect 2398 573 2432 679
rect 2556 573 2590 679
rect 2674 573 2708 679
rect 2832 573 2866 679
rect 2950 573 2984 679
rect 3108 573 3142 679
rect 3226 573 3260 679
rect 3384 573 3418 679
rect 3502 573 3536 679
rect 3660 573 3694 679
rect 3778 573 3812 679
rect 3936 573 3970 679
rect 4054 573 4088 679
rect 4212 573 4246 679
rect 4330 573 4364 679
rect 4488 573 4522 679
rect 4606 573 4640 679
rect 4764 573 4798 679
rect 4882 573 4916 679
rect 5040 573 5074 679
rect 5158 573 5192 679
rect 5316 573 5350 679
rect 252 489 320 523
rect 528 489 596 523
rect 804 489 872 523
rect 1080 489 1148 523
rect 1356 489 1424 523
rect 1632 489 1700 523
rect 1908 489 1976 523
rect 2184 489 2252 523
rect 2460 489 2528 523
rect 2736 489 2804 523
rect 3012 489 3080 523
rect 3288 489 3356 523
rect 3564 489 3632 523
rect 3840 489 3908 523
rect 4116 489 4184 523
rect 4392 489 4460 523
rect 4668 489 4736 523
rect 4944 489 5012 523
rect 5220 489 5288 523
rect 252 381 320 415
rect 528 381 596 415
rect 804 381 872 415
rect 1080 381 1148 415
rect 1356 381 1424 415
rect 1632 381 1700 415
rect 1908 381 1976 415
rect 2184 381 2252 415
rect 2460 381 2528 415
rect 2736 381 2804 415
rect 3012 381 3080 415
rect 3288 381 3356 415
rect 3564 381 3632 415
rect 3840 381 3908 415
rect 4116 381 4184 415
rect 4392 381 4460 415
rect 4668 381 4736 415
rect 4944 381 5012 415
rect 5220 381 5288 415
rect 190 225 224 331
rect 348 225 382 331
rect 466 225 500 331
rect 624 225 658 331
rect 742 225 776 331
rect 900 225 934 331
rect 1018 225 1052 331
rect 1176 225 1210 331
rect 1294 225 1328 331
rect 1452 225 1486 331
rect 1570 225 1604 331
rect 1728 225 1762 331
rect 1846 225 1880 331
rect 2004 225 2038 331
rect 2122 225 2156 331
rect 2280 225 2314 331
rect 2398 225 2432 331
rect 2556 225 2590 331
rect 2674 225 2708 331
rect 2832 225 2866 331
rect 2950 225 2984 331
rect 3108 225 3142 331
rect 3226 225 3260 331
rect 3384 225 3418 331
rect 3502 225 3536 331
rect 3660 225 3694 331
rect 3778 225 3812 331
rect 3936 225 3970 331
rect 4054 225 4088 331
rect 4212 225 4246 331
rect 4330 225 4364 331
rect 4488 225 4522 331
rect 4606 225 4640 331
rect 4764 225 4798 331
rect 4882 225 4916 331
rect 5040 225 5074 331
rect 5158 225 5192 331
rect 5316 225 5350 331
rect 252 141 320 175
rect 528 141 596 175
rect 804 141 872 175
rect 1080 141 1148 175
rect 1356 141 1424 175
rect 1632 141 1700 175
rect 1908 141 1976 175
rect 2184 141 2252 175
rect 2460 141 2528 175
rect 2736 141 2804 175
rect 3012 141 3080 175
rect 3288 141 3356 175
rect 3564 141 3632 175
rect 3840 141 3908 175
rect 4116 141 4184 175
rect 4392 141 4460 175
rect 4668 141 4736 175
rect 4944 141 5012 175
rect 5220 141 5288 175
rect 172 48 400 82
rect 448 48 676 82
rect 724 48 952 82
rect 1000 48 1228 82
rect 1276 48 1504 82
rect 1552 48 1780 82
rect 1828 48 2056 82
rect 2104 48 2332 82
rect 2380 48 2608 82
rect 2656 48 2884 82
rect 2932 48 3160 82
rect 3208 48 3436 82
rect 3484 48 3712 82
rect 3760 48 3988 82
rect 4036 48 4264 82
rect 4312 48 4540 82
rect 4588 48 4816 82
rect 4864 48 5092 82
rect 5140 48 5368 82
<< metal1 >>
rect 148 1998 5392 2010
rect 148 1964 172 1998
rect 400 1964 448 1998
rect 676 1964 724 1998
rect 952 1964 1000 1998
rect 1228 1964 1276 1998
rect 1504 1964 1552 1998
rect 1780 1964 1828 1998
rect 2056 1964 2104 1998
rect 2332 1964 2380 1998
rect 2608 1964 2656 1998
rect 2884 1964 2932 1998
rect 3160 1964 3208 1998
rect 3436 1964 3484 1998
rect 3712 1964 3760 1998
rect 3988 1964 4036 1998
rect 4264 1964 4312 1998
rect 4540 1964 4588 1998
rect 4816 1964 4864 1998
rect 5092 1964 5140 1998
rect 5368 1964 5392 1998
rect 148 1952 5392 1964
rect 240 1914 332 1920
rect 240 1880 252 1914
rect 320 1880 332 1914
rect 240 1874 332 1880
rect 516 1914 608 1920
rect 516 1880 528 1914
rect 596 1880 608 1914
rect 516 1874 608 1880
rect 792 1914 884 1920
rect 792 1880 804 1914
rect 872 1880 884 1914
rect 792 1874 884 1880
rect 1068 1914 1160 1920
rect 1068 1880 1080 1914
rect 1148 1880 1160 1914
rect 1068 1874 1160 1880
rect 1344 1914 1436 1920
rect 1344 1880 1356 1914
rect 1424 1880 1436 1914
rect 1344 1874 1436 1880
rect 1620 1914 1712 1920
rect 1620 1880 1632 1914
rect 1700 1880 1712 1914
rect 1620 1874 1712 1880
rect 1896 1914 1988 1920
rect 1896 1880 1908 1914
rect 1976 1880 1988 1914
rect 1896 1874 1988 1880
rect 2172 1914 2264 1920
rect 2172 1880 2184 1914
rect 2252 1880 2264 1914
rect 2172 1874 2264 1880
rect 2448 1914 2540 1920
rect 2448 1880 2460 1914
rect 2528 1880 2540 1914
rect 2448 1874 2540 1880
rect 2724 1914 2816 1920
rect 2724 1880 2736 1914
rect 2804 1880 2816 1914
rect 2724 1874 2816 1880
rect 3000 1914 3092 1920
rect 3000 1880 3012 1914
rect 3080 1880 3092 1914
rect 3000 1874 3092 1880
rect 3276 1914 3368 1920
rect 3276 1880 3288 1914
rect 3356 1880 3368 1914
rect 3276 1874 3368 1880
rect 3552 1914 3644 1920
rect 3552 1880 3564 1914
rect 3632 1880 3644 1914
rect 3552 1874 3644 1880
rect 3828 1914 3920 1920
rect 3828 1880 3840 1914
rect 3908 1880 3920 1914
rect 3828 1874 3920 1880
rect 4104 1914 4196 1920
rect 4104 1880 4116 1914
rect 4184 1880 4196 1914
rect 4104 1874 4196 1880
rect 4380 1914 4472 1920
rect 4380 1880 4392 1914
rect 4460 1880 4472 1914
rect 4380 1874 4472 1880
rect 4656 1914 4748 1920
rect 4656 1880 4668 1914
rect 4736 1880 4748 1914
rect 4656 1874 4748 1880
rect 4932 1914 5024 1920
rect 4932 1880 4944 1914
rect 5012 1880 5024 1914
rect 4932 1874 5024 1880
rect 5208 1914 5300 1920
rect 5208 1880 5220 1914
rect 5288 1880 5300 1914
rect 5208 1874 5300 1880
rect 184 1821 230 1833
rect 184 1645 190 1821
rect 224 1645 230 1821
rect 184 1633 230 1645
rect 269 1592 303 1874
rect 342 1821 388 1833
rect 342 1645 348 1821
rect 382 1645 388 1821
rect 342 1633 388 1645
rect 460 1821 506 1833
rect 460 1645 466 1821
rect 500 1645 506 1821
rect 460 1633 506 1645
rect 545 1592 579 1874
rect 618 1821 664 1833
rect 618 1645 624 1821
rect 658 1645 664 1821
rect 618 1633 664 1645
rect 736 1821 782 1833
rect 736 1645 742 1821
rect 776 1645 782 1821
rect 736 1633 782 1645
rect 821 1592 855 1874
rect 894 1821 940 1833
rect 894 1645 900 1821
rect 934 1645 940 1821
rect 894 1633 940 1645
rect 1012 1821 1058 1833
rect 1012 1645 1018 1821
rect 1052 1645 1058 1821
rect 1012 1633 1058 1645
rect 1097 1592 1131 1874
rect 1170 1821 1216 1833
rect 1170 1645 1176 1821
rect 1210 1645 1216 1821
rect 1170 1633 1216 1645
rect 1288 1821 1334 1833
rect 1288 1645 1294 1821
rect 1328 1645 1334 1821
rect 1288 1633 1334 1645
rect 1373 1592 1407 1874
rect 1446 1821 1492 1833
rect 1446 1645 1452 1821
rect 1486 1645 1492 1821
rect 1446 1633 1492 1645
rect 1564 1821 1610 1833
rect 1564 1645 1570 1821
rect 1604 1645 1610 1821
rect 1564 1633 1610 1645
rect 1649 1592 1683 1874
rect 1722 1821 1768 1833
rect 1722 1645 1728 1821
rect 1762 1645 1768 1821
rect 1722 1633 1768 1645
rect 1840 1821 1886 1833
rect 1840 1645 1846 1821
rect 1880 1645 1886 1821
rect 1840 1633 1886 1645
rect 1925 1592 1959 1874
rect 1998 1821 2044 1833
rect 1998 1645 2004 1821
rect 2038 1645 2044 1821
rect 1998 1633 2044 1645
rect 2116 1821 2162 1833
rect 2116 1645 2122 1821
rect 2156 1645 2162 1821
rect 2116 1633 2162 1645
rect 2201 1592 2235 1874
rect 2274 1821 2320 1833
rect 2274 1645 2280 1821
rect 2314 1645 2320 1821
rect 2274 1633 2320 1645
rect 2392 1821 2438 1833
rect 2392 1645 2398 1821
rect 2432 1645 2438 1821
rect 2392 1633 2438 1645
rect 2477 1592 2511 1874
rect 2550 1821 2596 1833
rect 2550 1645 2556 1821
rect 2590 1645 2596 1821
rect 2550 1633 2596 1645
rect 2668 1821 2714 1833
rect 2668 1645 2674 1821
rect 2708 1645 2714 1821
rect 2668 1633 2714 1645
rect 2753 1592 2787 1874
rect 2826 1821 2872 1833
rect 2826 1645 2832 1821
rect 2866 1645 2872 1821
rect 2826 1633 2872 1645
rect 2944 1821 2990 1833
rect 2944 1645 2950 1821
rect 2984 1645 2990 1821
rect 2944 1633 2990 1645
rect 3029 1592 3063 1874
rect 3102 1821 3148 1833
rect 3102 1645 3108 1821
rect 3142 1645 3148 1821
rect 3102 1633 3148 1645
rect 3220 1821 3266 1833
rect 3220 1645 3226 1821
rect 3260 1645 3266 1821
rect 3220 1633 3266 1645
rect 3305 1592 3339 1874
rect 3378 1821 3424 1833
rect 3378 1645 3384 1821
rect 3418 1645 3424 1821
rect 3378 1633 3424 1645
rect 3496 1821 3542 1833
rect 3496 1645 3502 1821
rect 3536 1645 3542 1821
rect 3496 1633 3542 1645
rect 3581 1592 3615 1874
rect 3654 1821 3700 1833
rect 3654 1645 3660 1821
rect 3694 1645 3700 1821
rect 3654 1633 3700 1645
rect 3772 1821 3818 1833
rect 3772 1645 3778 1821
rect 3812 1645 3818 1821
rect 3772 1633 3818 1645
rect 3857 1592 3891 1874
rect 3930 1821 3976 1833
rect 3930 1645 3936 1821
rect 3970 1645 3976 1821
rect 3930 1633 3976 1645
rect 4048 1821 4094 1833
rect 4048 1645 4054 1821
rect 4088 1645 4094 1821
rect 4048 1633 4094 1645
rect 4133 1592 4167 1874
rect 4206 1821 4252 1833
rect 4206 1645 4212 1821
rect 4246 1645 4252 1821
rect 4206 1633 4252 1645
rect 4324 1821 4370 1833
rect 4324 1645 4330 1821
rect 4364 1645 4370 1821
rect 4324 1633 4370 1645
rect 4409 1592 4443 1874
rect 4482 1821 4528 1833
rect 4482 1645 4488 1821
rect 4522 1645 4528 1821
rect 4482 1633 4528 1645
rect 4600 1821 4646 1833
rect 4600 1645 4606 1821
rect 4640 1645 4646 1821
rect 4600 1633 4646 1645
rect 4685 1592 4719 1874
rect 4758 1821 4804 1833
rect 4758 1645 4764 1821
rect 4798 1645 4804 1821
rect 4758 1633 4804 1645
rect 4876 1821 4922 1833
rect 4876 1645 4882 1821
rect 4916 1645 4922 1821
rect 4876 1633 4922 1645
rect 4961 1592 4995 1874
rect 5034 1821 5080 1833
rect 5034 1645 5040 1821
rect 5074 1645 5080 1821
rect 5034 1633 5080 1645
rect 5152 1821 5198 1833
rect 5152 1645 5158 1821
rect 5192 1645 5198 1821
rect 5152 1633 5198 1645
rect 5237 1592 5271 1874
rect 5310 1821 5356 1833
rect 5310 1645 5316 1821
rect 5350 1645 5356 1821
rect 5310 1633 5356 1645
rect 240 1586 332 1592
rect 240 1552 252 1586
rect 320 1552 332 1586
rect 240 1546 332 1552
rect 516 1586 608 1592
rect 516 1552 528 1586
rect 596 1552 608 1586
rect 516 1546 608 1552
rect 792 1586 884 1592
rect 792 1552 804 1586
rect 872 1552 884 1586
rect 792 1546 884 1552
rect 1068 1586 1160 1592
rect 1068 1552 1080 1586
rect 1148 1552 1160 1586
rect 1068 1546 1160 1552
rect 1344 1586 1436 1592
rect 1344 1552 1356 1586
rect 1424 1552 1436 1586
rect 1344 1546 1436 1552
rect 1620 1586 1712 1592
rect 1620 1552 1632 1586
rect 1700 1552 1712 1586
rect 1620 1546 1712 1552
rect 1896 1586 1988 1592
rect 1896 1552 1908 1586
rect 1976 1552 1988 1586
rect 1896 1546 1988 1552
rect 2172 1586 2264 1592
rect 2172 1552 2184 1586
rect 2252 1552 2264 1586
rect 2172 1546 2264 1552
rect 2448 1586 2540 1592
rect 2448 1552 2460 1586
rect 2528 1552 2540 1586
rect 2448 1546 2540 1552
rect 2724 1586 2816 1592
rect 2724 1552 2736 1586
rect 2804 1552 2816 1586
rect 2724 1546 2816 1552
rect 3000 1586 3092 1592
rect 3000 1552 3012 1586
rect 3080 1552 3092 1586
rect 3000 1546 3092 1552
rect 3276 1586 3368 1592
rect 3276 1552 3288 1586
rect 3356 1552 3368 1586
rect 3276 1546 3368 1552
rect 3552 1586 3644 1592
rect 3552 1552 3564 1586
rect 3632 1552 3644 1586
rect 3552 1546 3644 1552
rect 3828 1586 3920 1592
rect 3828 1552 3840 1586
rect 3908 1552 3920 1586
rect 3828 1546 3920 1552
rect 4104 1586 4196 1592
rect 4104 1552 4116 1586
rect 4184 1552 4196 1586
rect 4104 1546 4196 1552
rect 4380 1586 4472 1592
rect 4380 1552 4392 1586
rect 4460 1552 4472 1586
rect 4380 1546 4472 1552
rect 4656 1586 4748 1592
rect 4656 1552 4668 1586
rect 4736 1552 4748 1586
rect 4656 1546 4748 1552
rect 4932 1586 5024 1592
rect 4932 1552 4944 1586
rect 5012 1552 5024 1586
rect 4932 1546 5024 1552
rect 5208 1586 5300 1592
rect 5208 1552 5220 1586
rect 5288 1552 5300 1586
rect 5208 1546 5300 1552
rect 240 1478 332 1484
rect 240 1444 252 1478
rect 320 1444 332 1478
rect 240 1438 332 1444
rect 516 1478 608 1484
rect 516 1444 528 1478
rect 596 1444 608 1478
rect 516 1438 608 1444
rect 792 1478 884 1484
rect 792 1444 804 1478
rect 872 1444 884 1478
rect 792 1438 884 1444
rect 1068 1478 1160 1484
rect 1068 1444 1080 1478
rect 1148 1444 1160 1478
rect 1068 1438 1160 1444
rect 1344 1478 1436 1484
rect 1344 1444 1356 1478
rect 1424 1444 1436 1478
rect 1344 1438 1436 1444
rect 1620 1478 1712 1484
rect 1620 1444 1632 1478
rect 1700 1444 1712 1478
rect 1620 1438 1712 1444
rect 1896 1478 1988 1484
rect 1896 1444 1908 1478
rect 1976 1444 1988 1478
rect 1896 1438 1988 1444
rect 2172 1478 2264 1484
rect 2172 1444 2184 1478
rect 2252 1444 2264 1478
rect 2172 1438 2264 1444
rect 2448 1478 2540 1484
rect 2448 1444 2460 1478
rect 2528 1444 2540 1478
rect 2448 1438 2540 1444
rect 2724 1478 2816 1484
rect 2724 1444 2736 1478
rect 2804 1444 2816 1478
rect 2724 1438 2816 1444
rect 3000 1478 3092 1484
rect 3000 1444 3012 1478
rect 3080 1444 3092 1478
rect 3000 1438 3092 1444
rect 3276 1478 3368 1484
rect 3276 1444 3288 1478
rect 3356 1444 3368 1478
rect 3276 1438 3368 1444
rect 3552 1478 3644 1484
rect 3552 1444 3564 1478
rect 3632 1444 3644 1478
rect 3552 1438 3644 1444
rect 3828 1478 3920 1484
rect 3828 1444 3840 1478
rect 3908 1444 3920 1478
rect 3828 1438 3920 1444
rect 4104 1478 4196 1484
rect 4104 1444 4116 1478
rect 4184 1444 4196 1478
rect 4104 1438 4196 1444
rect 4380 1478 4472 1484
rect 4380 1444 4392 1478
rect 4460 1444 4472 1478
rect 4380 1438 4472 1444
rect 4656 1478 4748 1484
rect 4656 1444 4668 1478
rect 4736 1444 4748 1478
rect 4656 1438 4748 1444
rect 4932 1478 5024 1484
rect 4932 1444 4944 1478
rect 5012 1444 5024 1478
rect 4932 1438 5024 1444
rect 5208 1478 5300 1484
rect 5208 1444 5220 1478
rect 5288 1444 5300 1478
rect 5208 1438 5300 1444
rect 184 1385 230 1397
rect 184 1209 190 1385
rect 224 1209 230 1385
rect 184 1197 230 1209
rect 269 1156 303 1438
rect 342 1385 388 1397
rect 342 1209 348 1385
rect 382 1209 388 1385
rect 342 1197 388 1209
rect 460 1385 506 1397
rect 460 1209 466 1385
rect 500 1209 506 1385
rect 460 1197 506 1209
rect 545 1156 579 1438
rect 618 1385 664 1397
rect 618 1209 624 1385
rect 658 1209 664 1385
rect 618 1197 664 1209
rect 736 1385 782 1397
rect 736 1209 742 1385
rect 776 1209 782 1385
rect 736 1197 782 1209
rect 821 1156 855 1438
rect 894 1385 940 1397
rect 894 1209 900 1385
rect 934 1209 940 1385
rect 894 1197 940 1209
rect 1012 1385 1058 1397
rect 1012 1209 1018 1385
rect 1052 1209 1058 1385
rect 1012 1197 1058 1209
rect 1097 1156 1131 1438
rect 1170 1385 1216 1397
rect 1170 1209 1176 1385
rect 1210 1209 1216 1385
rect 1170 1197 1216 1209
rect 1288 1385 1334 1397
rect 1288 1209 1294 1385
rect 1328 1209 1334 1385
rect 1288 1197 1334 1209
rect 1373 1156 1407 1438
rect 1446 1385 1492 1397
rect 1446 1209 1452 1385
rect 1486 1209 1492 1385
rect 1446 1197 1492 1209
rect 1564 1385 1610 1397
rect 1564 1209 1570 1385
rect 1604 1209 1610 1385
rect 1564 1197 1610 1209
rect 1649 1156 1683 1438
rect 1722 1385 1768 1397
rect 1722 1209 1728 1385
rect 1762 1209 1768 1385
rect 1722 1197 1768 1209
rect 1840 1385 1886 1397
rect 1840 1209 1846 1385
rect 1880 1209 1886 1385
rect 1840 1197 1886 1209
rect 1925 1156 1959 1438
rect 1998 1385 2044 1397
rect 1998 1209 2004 1385
rect 2038 1209 2044 1385
rect 1998 1197 2044 1209
rect 2116 1385 2162 1397
rect 2116 1209 2122 1385
rect 2156 1209 2162 1385
rect 2116 1197 2162 1209
rect 2201 1156 2235 1438
rect 2274 1385 2320 1397
rect 2274 1209 2280 1385
rect 2314 1209 2320 1385
rect 2274 1197 2320 1209
rect 2392 1385 2438 1397
rect 2392 1209 2398 1385
rect 2432 1209 2438 1385
rect 2392 1197 2438 1209
rect 2477 1156 2511 1438
rect 2550 1385 2596 1397
rect 2550 1209 2556 1385
rect 2590 1209 2596 1385
rect 2550 1197 2596 1209
rect 2668 1385 2714 1397
rect 2668 1209 2674 1385
rect 2708 1209 2714 1385
rect 2668 1197 2714 1209
rect 2753 1156 2787 1438
rect 2826 1385 2872 1397
rect 2826 1209 2832 1385
rect 2866 1209 2872 1385
rect 2826 1197 2872 1209
rect 2944 1385 2990 1397
rect 2944 1209 2950 1385
rect 2984 1209 2990 1385
rect 2944 1197 2990 1209
rect 3029 1156 3063 1438
rect 3102 1385 3148 1397
rect 3102 1209 3108 1385
rect 3142 1209 3148 1385
rect 3102 1197 3148 1209
rect 3220 1385 3266 1397
rect 3220 1209 3226 1385
rect 3260 1209 3266 1385
rect 3220 1197 3266 1209
rect 3305 1156 3339 1438
rect 3378 1385 3424 1397
rect 3378 1209 3384 1385
rect 3418 1209 3424 1385
rect 3378 1197 3424 1209
rect 3496 1385 3542 1397
rect 3496 1209 3502 1385
rect 3536 1209 3542 1385
rect 3496 1197 3542 1209
rect 3581 1156 3615 1438
rect 3654 1385 3700 1397
rect 3654 1209 3660 1385
rect 3694 1209 3700 1385
rect 3654 1197 3700 1209
rect 3772 1385 3818 1397
rect 3772 1209 3778 1385
rect 3812 1209 3818 1385
rect 3772 1197 3818 1209
rect 3857 1156 3891 1438
rect 3930 1385 3976 1397
rect 3930 1209 3936 1385
rect 3970 1209 3976 1385
rect 3930 1197 3976 1209
rect 4048 1385 4094 1397
rect 4048 1209 4054 1385
rect 4088 1209 4094 1385
rect 4048 1197 4094 1209
rect 4133 1156 4167 1438
rect 4206 1385 4252 1397
rect 4206 1209 4212 1385
rect 4246 1209 4252 1385
rect 4206 1197 4252 1209
rect 4324 1385 4370 1397
rect 4324 1209 4330 1385
rect 4364 1209 4370 1385
rect 4324 1197 4370 1209
rect 4409 1156 4443 1438
rect 4482 1385 4528 1397
rect 4482 1209 4488 1385
rect 4522 1209 4528 1385
rect 4482 1197 4528 1209
rect 4600 1385 4646 1397
rect 4600 1209 4606 1385
rect 4640 1209 4646 1385
rect 4600 1197 4646 1209
rect 4685 1156 4719 1438
rect 4758 1385 4804 1397
rect 4758 1209 4764 1385
rect 4798 1209 4804 1385
rect 4758 1197 4804 1209
rect 4876 1385 4922 1397
rect 4876 1209 4882 1385
rect 4916 1209 4922 1385
rect 4876 1197 4922 1209
rect 4961 1156 4995 1438
rect 5034 1385 5080 1397
rect 5034 1209 5040 1385
rect 5074 1209 5080 1385
rect 5034 1197 5080 1209
rect 5152 1385 5198 1397
rect 5152 1209 5158 1385
rect 5192 1209 5198 1385
rect 5152 1197 5198 1209
rect 5237 1156 5271 1438
rect 5310 1385 5356 1397
rect 5310 1209 5316 1385
rect 5350 1209 5356 1385
rect 5310 1197 5356 1209
rect 240 1150 332 1156
rect 240 1116 252 1150
rect 320 1116 332 1150
rect 240 1110 332 1116
rect 516 1150 608 1156
rect 516 1116 528 1150
rect 596 1116 608 1150
rect 516 1110 608 1116
rect 792 1150 884 1156
rect 792 1116 804 1150
rect 872 1116 884 1150
rect 792 1110 884 1116
rect 1068 1150 1160 1156
rect 1068 1116 1080 1150
rect 1148 1116 1160 1150
rect 1068 1110 1160 1116
rect 1344 1150 1436 1156
rect 1344 1116 1356 1150
rect 1424 1116 1436 1150
rect 1344 1110 1436 1116
rect 1620 1150 1712 1156
rect 1620 1116 1632 1150
rect 1700 1116 1712 1150
rect 1620 1110 1712 1116
rect 1896 1150 1988 1156
rect 1896 1116 1908 1150
rect 1976 1116 1988 1150
rect 1896 1110 1988 1116
rect 2172 1150 2264 1156
rect 2172 1116 2184 1150
rect 2252 1116 2264 1150
rect 2172 1110 2264 1116
rect 2448 1150 2540 1156
rect 2448 1116 2460 1150
rect 2528 1116 2540 1150
rect 2448 1110 2540 1116
rect 2724 1150 2816 1156
rect 2724 1116 2736 1150
rect 2804 1116 2816 1150
rect 2724 1110 2816 1116
rect 3000 1150 3092 1156
rect 3000 1116 3012 1150
rect 3080 1116 3092 1150
rect 3000 1110 3092 1116
rect 3276 1150 3368 1156
rect 3276 1116 3288 1150
rect 3356 1116 3368 1150
rect 3276 1110 3368 1116
rect 3552 1150 3644 1156
rect 3552 1116 3564 1150
rect 3632 1116 3644 1150
rect 3552 1110 3644 1116
rect 3828 1150 3920 1156
rect 3828 1116 3840 1150
rect 3908 1116 3920 1150
rect 3828 1110 3920 1116
rect 4104 1150 4196 1156
rect 4104 1116 4116 1150
rect 4184 1116 4196 1150
rect 4104 1110 4196 1116
rect 4380 1150 4472 1156
rect 4380 1116 4392 1150
rect 4460 1116 4472 1150
rect 4380 1110 4472 1116
rect 4656 1150 4748 1156
rect 4656 1116 4668 1150
rect 4736 1116 4748 1150
rect 4656 1110 4748 1116
rect 4932 1150 5024 1156
rect 4932 1116 4944 1150
rect 5012 1116 5024 1150
rect 4932 1110 5024 1116
rect 5208 1150 5300 1156
rect 5208 1116 5220 1150
rect 5288 1116 5300 1150
rect 5208 1110 5300 1116
rect 240 763 332 769
rect 240 729 252 763
rect 320 729 332 763
rect 240 723 332 729
rect 516 763 608 769
rect 516 729 528 763
rect 596 729 608 763
rect 516 723 608 729
rect 792 763 884 769
rect 792 729 804 763
rect 872 729 884 763
rect 792 723 884 729
rect 1068 763 1160 769
rect 1068 729 1080 763
rect 1148 729 1160 763
rect 1068 723 1160 729
rect 1344 763 1436 769
rect 1344 729 1356 763
rect 1424 729 1436 763
rect 1344 723 1436 729
rect 1620 763 1712 769
rect 1620 729 1632 763
rect 1700 729 1712 763
rect 1620 723 1712 729
rect 1896 763 1988 769
rect 1896 729 1908 763
rect 1976 729 1988 763
rect 1896 723 1988 729
rect 2172 763 2264 769
rect 2172 729 2184 763
rect 2252 729 2264 763
rect 2172 723 2264 729
rect 2448 763 2540 769
rect 2448 729 2460 763
rect 2528 729 2540 763
rect 2448 723 2540 729
rect 2724 763 2816 769
rect 2724 729 2736 763
rect 2804 729 2816 763
rect 2724 723 2816 729
rect 3000 763 3092 769
rect 3000 729 3012 763
rect 3080 729 3092 763
rect 3000 723 3092 729
rect 3276 763 3368 769
rect 3276 729 3288 763
rect 3356 729 3368 763
rect 3276 723 3368 729
rect 3552 763 3644 769
rect 3552 729 3564 763
rect 3632 729 3644 763
rect 3552 723 3644 729
rect 3828 763 3920 769
rect 3828 729 3840 763
rect 3908 729 3920 763
rect 3828 723 3920 729
rect 4104 763 4196 769
rect 4104 729 4116 763
rect 4184 729 4196 763
rect 4104 723 4196 729
rect 4380 763 4472 769
rect 4380 729 4392 763
rect 4460 729 4472 763
rect 4380 723 4472 729
rect 4656 763 4748 769
rect 4656 729 4668 763
rect 4736 729 4748 763
rect 4656 723 4748 729
rect 4932 763 5024 769
rect 4932 729 4944 763
rect 5012 729 5024 763
rect 4932 723 5024 729
rect 5208 763 5300 769
rect 5208 729 5220 763
rect 5288 729 5300 763
rect 5208 723 5300 729
rect 184 679 230 691
rect 184 573 190 679
rect 224 573 230 679
rect 184 561 230 573
rect 269 529 303 723
rect 342 679 388 691
rect 342 573 348 679
rect 382 573 388 679
rect 342 561 388 573
rect 460 679 506 691
rect 460 573 466 679
rect 500 573 506 679
rect 460 561 506 573
rect 545 529 579 723
rect 618 679 664 691
rect 618 573 624 679
rect 658 573 664 679
rect 618 561 664 573
rect 736 679 782 691
rect 736 573 742 679
rect 776 573 782 679
rect 736 561 782 573
rect 821 529 855 723
rect 894 679 940 691
rect 894 573 900 679
rect 934 573 940 679
rect 894 561 940 573
rect 1012 679 1058 691
rect 1012 573 1018 679
rect 1052 573 1058 679
rect 1012 561 1058 573
rect 1097 529 1131 723
rect 1170 679 1216 691
rect 1170 573 1176 679
rect 1210 573 1216 679
rect 1170 561 1216 573
rect 1288 679 1334 691
rect 1288 573 1294 679
rect 1328 573 1334 679
rect 1288 561 1334 573
rect 1373 529 1407 723
rect 1446 679 1492 691
rect 1446 573 1452 679
rect 1486 573 1492 679
rect 1446 561 1492 573
rect 1564 679 1610 691
rect 1564 573 1570 679
rect 1604 573 1610 679
rect 1564 561 1610 573
rect 1649 529 1683 723
rect 1722 679 1768 691
rect 1722 573 1728 679
rect 1762 573 1768 679
rect 1722 561 1768 573
rect 1840 679 1886 691
rect 1840 573 1846 679
rect 1880 573 1886 679
rect 1840 561 1886 573
rect 1925 529 1959 723
rect 1998 679 2044 691
rect 1998 573 2004 679
rect 2038 573 2044 679
rect 1998 561 2044 573
rect 2116 679 2162 691
rect 2116 573 2122 679
rect 2156 573 2162 679
rect 2116 561 2162 573
rect 2201 529 2235 723
rect 2274 679 2320 691
rect 2274 573 2280 679
rect 2314 573 2320 679
rect 2274 561 2320 573
rect 2392 679 2438 691
rect 2392 573 2398 679
rect 2432 573 2438 679
rect 2392 561 2438 573
rect 2477 529 2511 723
rect 2550 679 2596 691
rect 2550 573 2556 679
rect 2590 573 2596 679
rect 2550 561 2596 573
rect 2668 679 2714 691
rect 2668 573 2674 679
rect 2708 573 2714 679
rect 2668 561 2714 573
rect 2753 529 2787 723
rect 2826 679 2872 691
rect 2826 573 2832 679
rect 2866 573 2872 679
rect 2826 561 2872 573
rect 2944 679 2990 691
rect 2944 573 2950 679
rect 2984 573 2990 679
rect 2944 561 2990 573
rect 3029 529 3063 723
rect 3102 679 3148 691
rect 3102 573 3108 679
rect 3142 573 3148 679
rect 3102 561 3148 573
rect 3220 679 3266 691
rect 3220 573 3226 679
rect 3260 573 3266 679
rect 3220 561 3266 573
rect 3305 529 3339 723
rect 3378 679 3424 691
rect 3378 573 3384 679
rect 3418 573 3424 679
rect 3378 561 3424 573
rect 3496 679 3542 691
rect 3496 573 3502 679
rect 3536 573 3542 679
rect 3496 561 3542 573
rect 3581 529 3615 723
rect 3654 679 3700 691
rect 3654 573 3660 679
rect 3694 573 3700 679
rect 3654 561 3700 573
rect 3772 679 3818 691
rect 3772 573 3778 679
rect 3812 573 3818 679
rect 3772 561 3818 573
rect 3857 529 3891 723
rect 3930 679 3976 691
rect 3930 573 3936 679
rect 3970 573 3976 679
rect 3930 561 3976 573
rect 4048 679 4094 691
rect 4048 573 4054 679
rect 4088 573 4094 679
rect 4048 561 4094 573
rect 4133 529 4167 723
rect 4206 679 4252 691
rect 4206 573 4212 679
rect 4246 573 4252 679
rect 4206 561 4252 573
rect 4324 679 4370 691
rect 4324 573 4330 679
rect 4364 573 4370 679
rect 4324 561 4370 573
rect 4409 529 4443 723
rect 4482 679 4528 691
rect 4482 573 4488 679
rect 4522 573 4528 679
rect 4482 561 4528 573
rect 4600 679 4646 691
rect 4600 573 4606 679
rect 4640 573 4646 679
rect 4600 561 4646 573
rect 4685 529 4719 723
rect 4758 679 4804 691
rect 4758 573 4764 679
rect 4798 573 4804 679
rect 4758 561 4804 573
rect 4876 679 4922 691
rect 4876 573 4882 679
rect 4916 573 4922 679
rect 4876 561 4922 573
rect 4961 529 4995 723
rect 5034 679 5080 691
rect 5034 573 5040 679
rect 5074 573 5080 679
rect 5034 561 5080 573
rect 5152 679 5198 691
rect 5152 573 5158 679
rect 5192 573 5198 679
rect 5152 561 5198 573
rect 5237 529 5271 723
rect 5310 679 5356 691
rect 5310 573 5316 679
rect 5350 573 5356 679
rect 5310 561 5356 573
rect 240 523 332 529
rect 240 489 252 523
rect 320 489 332 523
rect 240 483 332 489
rect 516 523 608 529
rect 516 489 528 523
rect 596 489 608 523
rect 516 483 608 489
rect 792 523 884 529
rect 792 489 804 523
rect 872 489 884 523
rect 792 483 884 489
rect 1068 523 1160 529
rect 1068 489 1080 523
rect 1148 489 1160 523
rect 1068 483 1160 489
rect 1344 523 1436 529
rect 1344 489 1356 523
rect 1424 489 1436 523
rect 1344 483 1436 489
rect 1620 523 1712 529
rect 1620 489 1632 523
rect 1700 489 1712 523
rect 1620 483 1712 489
rect 1896 523 1988 529
rect 1896 489 1908 523
rect 1976 489 1988 523
rect 1896 483 1988 489
rect 2172 523 2264 529
rect 2172 489 2184 523
rect 2252 489 2264 523
rect 2172 483 2264 489
rect 2448 523 2540 529
rect 2448 489 2460 523
rect 2528 489 2540 523
rect 2448 483 2540 489
rect 2724 523 2816 529
rect 2724 489 2736 523
rect 2804 489 2816 523
rect 2724 483 2816 489
rect 3000 523 3092 529
rect 3000 489 3012 523
rect 3080 489 3092 523
rect 3000 483 3092 489
rect 3276 523 3368 529
rect 3276 489 3288 523
rect 3356 489 3368 523
rect 3276 483 3368 489
rect 3552 523 3644 529
rect 3552 489 3564 523
rect 3632 489 3644 523
rect 3552 483 3644 489
rect 3828 523 3920 529
rect 3828 489 3840 523
rect 3908 489 3920 523
rect 3828 483 3920 489
rect 4104 523 4196 529
rect 4104 489 4116 523
rect 4184 489 4196 523
rect 4104 483 4196 489
rect 4380 523 4472 529
rect 4380 489 4392 523
rect 4460 489 4472 523
rect 4380 483 4472 489
rect 4656 523 4748 529
rect 4656 489 4668 523
rect 4736 489 4748 523
rect 4656 483 4748 489
rect 4932 523 5024 529
rect 4932 489 4944 523
rect 5012 489 5024 523
rect 4932 483 5024 489
rect 5208 523 5300 529
rect 5208 489 5220 523
rect 5288 489 5300 523
rect 5208 483 5300 489
rect 240 415 332 421
rect 240 381 252 415
rect 320 381 332 415
rect 240 375 332 381
rect 516 415 608 421
rect 516 381 528 415
rect 596 381 608 415
rect 516 375 608 381
rect 792 415 884 421
rect 792 381 804 415
rect 872 381 884 415
rect 792 375 884 381
rect 1068 415 1160 421
rect 1068 381 1080 415
rect 1148 381 1160 415
rect 1068 375 1160 381
rect 1344 415 1436 421
rect 1344 381 1356 415
rect 1424 381 1436 415
rect 1344 375 1436 381
rect 1620 415 1712 421
rect 1620 381 1632 415
rect 1700 381 1712 415
rect 1620 375 1712 381
rect 1896 415 1988 421
rect 1896 381 1908 415
rect 1976 381 1988 415
rect 1896 375 1988 381
rect 2172 415 2264 421
rect 2172 381 2184 415
rect 2252 381 2264 415
rect 2172 375 2264 381
rect 2448 415 2540 421
rect 2448 381 2460 415
rect 2528 381 2540 415
rect 2448 375 2540 381
rect 2724 415 2816 421
rect 2724 381 2736 415
rect 2804 381 2816 415
rect 2724 375 2816 381
rect 3000 415 3092 421
rect 3000 381 3012 415
rect 3080 381 3092 415
rect 3000 375 3092 381
rect 3276 415 3368 421
rect 3276 381 3288 415
rect 3356 381 3368 415
rect 3276 375 3368 381
rect 3552 415 3644 421
rect 3552 381 3564 415
rect 3632 381 3644 415
rect 3552 375 3644 381
rect 3828 415 3920 421
rect 3828 381 3840 415
rect 3908 381 3920 415
rect 3828 375 3920 381
rect 4104 415 4196 421
rect 4104 381 4116 415
rect 4184 381 4196 415
rect 4104 375 4196 381
rect 4380 415 4472 421
rect 4380 381 4392 415
rect 4460 381 4472 415
rect 4380 375 4472 381
rect 4656 415 4748 421
rect 4656 381 4668 415
rect 4736 381 4748 415
rect 4656 375 4748 381
rect 4932 415 5024 421
rect 4932 381 4944 415
rect 5012 381 5024 415
rect 4932 375 5024 381
rect 5208 415 5300 421
rect 5208 381 5220 415
rect 5288 381 5300 415
rect 5208 375 5300 381
rect 184 331 230 343
rect 184 225 190 331
rect 224 225 230 331
rect 184 213 230 225
rect 269 181 303 375
rect 342 331 388 343
rect 342 225 348 331
rect 382 225 388 331
rect 342 213 388 225
rect 460 331 506 343
rect 460 225 466 331
rect 500 225 506 331
rect 460 213 506 225
rect 545 181 579 375
rect 618 331 664 343
rect 618 225 624 331
rect 658 225 664 331
rect 618 213 664 225
rect 736 331 782 343
rect 736 225 742 331
rect 776 225 782 331
rect 736 213 782 225
rect 821 181 855 375
rect 894 331 940 343
rect 894 225 900 331
rect 934 225 940 331
rect 894 213 940 225
rect 1012 331 1058 343
rect 1012 225 1018 331
rect 1052 225 1058 331
rect 1012 213 1058 225
rect 1097 181 1131 375
rect 1170 331 1216 343
rect 1170 225 1176 331
rect 1210 225 1216 331
rect 1170 213 1216 225
rect 1288 331 1334 343
rect 1288 225 1294 331
rect 1328 225 1334 331
rect 1288 213 1334 225
rect 1373 181 1407 375
rect 1446 331 1492 343
rect 1446 225 1452 331
rect 1486 225 1492 331
rect 1446 213 1492 225
rect 1564 331 1610 343
rect 1564 225 1570 331
rect 1604 225 1610 331
rect 1564 213 1610 225
rect 1649 181 1683 375
rect 1722 331 1768 343
rect 1722 225 1728 331
rect 1762 225 1768 331
rect 1722 213 1768 225
rect 1840 331 1886 343
rect 1840 225 1846 331
rect 1880 225 1886 331
rect 1840 213 1886 225
rect 1925 181 1959 375
rect 1998 331 2044 343
rect 1998 225 2004 331
rect 2038 225 2044 331
rect 1998 213 2044 225
rect 2116 331 2162 343
rect 2116 225 2122 331
rect 2156 225 2162 331
rect 2116 213 2162 225
rect 2201 181 2235 375
rect 2274 331 2320 343
rect 2274 225 2280 331
rect 2314 225 2320 331
rect 2274 213 2320 225
rect 2392 331 2438 343
rect 2392 225 2398 331
rect 2432 225 2438 331
rect 2392 213 2438 225
rect 2477 181 2511 375
rect 2550 331 2596 343
rect 2550 225 2556 331
rect 2590 225 2596 331
rect 2550 213 2596 225
rect 2668 331 2714 343
rect 2668 225 2674 331
rect 2708 225 2714 331
rect 2668 213 2714 225
rect 2753 181 2787 375
rect 2826 331 2872 343
rect 2826 225 2832 331
rect 2866 225 2872 331
rect 2826 213 2872 225
rect 2944 331 2990 343
rect 2944 225 2950 331
rect 2984 225 2990 331
rect 2944 213 2990 225
rect 3029 181 3063 375
rect 3102 331 3148 343
rect 3102 225 3108 331
rect 3142 225 3148 331
rect 3102 213 3148 225
rect 3220 331 3266 343
rect 3220 225 3226 331
rect 3260 225 3266 331
rect 3220 213 3266 225
rect 3305 181 3339 375
rect 3378 331 3424 343
rect 3378 225 3384 331
rect 3418 225 3424 331
rect 3378 213 3424 225
rect 3496 331 3542 343
rect 3496 225 3502 331
rect 3536 225 3542 331
rect 3496 213 3542 225
rect 3581 181 3615 375
rect 3654 331 3700 343
rect 3654 225 3660 331
rect 3694 225 3700 331
rect 3654 213 3700 225
rect 3772 331 3818 343
rect 3772 225 3778 331
rect 3812 225 3818 331
rect 3772 213 3818 225
rect 3857 181 3891 375
rect 3930 331 3976 343
rect 3930 225 3936 331
rect 3970 225 3976 331
rect 3930 213 3976 225
rect 4048 331 4094 343
rect 4048 225 4054 331
rect 4088 225 4094 331
rect 4048 213 4094 225
rect 4133 181 4167 375
rect 4206 331 4252 343
rect 4206 225 4212 331
rect 4246 225 4252 331
rect 4206 213 4252 225
rect 4324 331 4370 343
rect 4324 225 4330 331
rect 4364 225 4370 331
rect 4324 213 4370 225
rect 4409 181 4443 375
rect 4482 331 4528 343
rect 4482 225 4488 331
rect 4522 225 4528 331
rect 4482 213 4528 225
rect 4600 331 4646 343
rect 4600 225 4606 331
rect 4640 225 4646 331
rect 4600 213 4646 225
rect 4685 181 4719 375
rect 4758 331 4804 343
rect 4758 225 4764 331
rect 4798 225 4804 331
rect 4758 213 4804 225
rect 4876 331 4922 343
rect 4876 225 4882 331
rect 4916 225 4922 331
rect 4876 213 4922 225
rect 4961 181 4995 375
rect 5034 331 5080 343
rect 5034 225 5040 331
rect 5074 225 5080 331
rect 5034 213 5080 225
rect 5152 331 5198 343
rect 5152 225 5158 331
rect 5192 225 5198 331
rect 5152 213 5198 225
rect 5237 181 5271 375
rect 5310 331 5356 343
rect 5310 225 5316 331
rect 5350 225 5356 331
rect 5310 213 5356 225
rect 240 175 332 181
rect 240 141 252 175
rect 320 141 332 175
rect 240 135 332 141
rect 516 175 608 181
rect 516 141 528 175
rect 596 141 608 175
rect 516 135 608 141
rect 792 175 884 181
rect 792 141 804 175
rect 872 141 884 175
rect 792 135 884 141
rect 1068 175 1160 181
rect 1068 141 1080 175
rect 1148 141 1160 175
rect 1068 135 1160 141
rect 1344 175 1436 181
rect 1344 141 1356 175
rect 1424 141 1436 175
rect 1344 135 1436 141
rect 1620 175 1712 181
rect 1620 141 1632 175
rect 1700 141 1712 175
rect 1620 135 1712 141
rect 1896 175 1988 181
rect 1896 141 1908 175
rect 1976 141 1988 175
rect 1896 135 1988 141
rect 2172 175 2264 181
rect 2172 141 2184 175
rect 2252 141 2264 175
rect 2172 135 2264 141
rect 2448 175 2540 181
rect 2448 141 2460 175
rect 2528 141 2540 175
rect 2448 135 2540 141
rect 2724 175 2816 181
rect 2724 141 2736 175
rect 2804 141 2816 175
rect 2724 135 2816 141
rect 3000 175 3092 181
rect 3000 141 3012 175
rect 3080 141 3092 175
rect 3000 135 3092 141
rect 3276 175 3368 181
rect 3276 141 3288 175
rect 3356 141 3368 175
rect 3276 135 3368 141
rect 3552 175 3644 181
rect 3552 141 3564 175
rect 3632 141 3644 175
rect 3552 135 3644 141
rect 3828 175 3920 181
rect 3828 141 3840 175
rect 3908 141 3920 175
rect 3828 135 3920 141
rect 4104 175 4196 181
rect 4104 141 4116 175
rect 4184 141 4196 175
rect 4104 135 4196 141
rect 4380 175 4472 181
rect 4380 141 4392 175
rect 4460 141 4472 175
rect 4380 135 4472 141
rect 4656 175 4748 181
rect 4656 141 4668 175
rect 4736 141 4748 175
rect 4656 135 4748 141
rect 4932 175 5024 181
rect 4932 141 4944 175
rect 5012 141 5024 175
rect 4932 135 5024 141
rect 5208 175 5300 181
rect 5208 141 5220 175
rect 5288 141 5300 175
rect 5208 135 5300 141
rect 148 82 5392 94
rect 148 48 172 82
rect 400 48 448 82
rect 676 48 724 82
rect 952 48 1000 82
rect 1228 48 1276 82
rect 1504 48 1552 82
rect 1780 48 1828 82
rect 2056 48 2104 82
rect 2332 48 2380 82
rect 2608 48 2656 82
rect 2884 48 2932 82
rect 3160 48 3208 82
rect 3436 48 3484 82
rect 3712 48 3760 82
rect 3988 48 4036 82
rect 4264 48 4312 82
rect 4540 48 4588 82
rect 4816 48 4864 82
rect 5092 48 5140 82
rect 5368 48 5392 82
rect 148 36 5392 48
<< labels >>
flabel metal1 148 1952 5392 2010 0 FreeSans 256 0 0 0 VDD
port 1 nsew power bidirectional
flabel metal1 148 36 5392 94 0 FreeSans 256 0 0 0 VSS
port 0 nsew ground bidirectional
<< end >>
