magic
tech sky130A
magscale 1 2
timestamp 1748318706
<< metal1 >>
rect 148 1168 2524 1226
rect 281 141 315 1130
rect 581 141 615 1130
rect 2472 209 2506 1053
rect 148 36 2524 94
use transistor_pair_bus_8  transistor_pair_bus_8_0
timestamp 1748299149
transform 1 0 60 0 1 0
box -60 0 2636 1292
use xor2_raw  xor2_raw_0
timestamp 1748318706
transform 1 0 0 0 1 0
box 148 36 2524 1226
<< labels >>
flabel metal1 281 141 315 1130 0 FreeSans 256 0 0 0 A
port 2 nsew signal input
flabel metal1 581 141 615 1130 0 FreeSans 256 0 0 0 B
port 3 nsew signal input
flabel metal1 2472 209 2506 1053 0 FreeSans 128 0 0 0 OUT
port 4 nsew signal output
flabel metal1 148 36 2524 94 0 FreeSans 256 0 0 0 VSS
port 0 nsew ground bidirectional
flabel metal1 148 1168 2524 1226 0 FreeSans 256 0 0 0 VDD
port 1 nsew power bidirectional
<< end >>
