magic
tech sky130A
magscale 1 2
timestamp 1748338064
<< metal1 >>
rect 4807 20378 4813 20430
rect 4865 20378 4871 20430
rect 7503 20378 7509 20430
rect 7561 20378 7567 20430
rect 10199 20378 10205 20430
rect 10257 20378 10263 20430
rect 12595 20384 12601 20436
rect 12653 20384 12659 20436
rect 12895 20378 12901 20430
rect 12953 20378 12959 20430
rect 5899 15862 5951 15868
rect 13776 15862 13828 15868
rect 5951 15819 13776 15853
rect 5899 15804 5951 15810
rect 13776 15804 13828 15810
rect 6175 15785 6227 15791
rect 14473 15785 14525 15791
rect 6227 15742 14473 15776
rect 6175 15727 6227 15733
rect 14473 15727 14525 15733
rect 6451 15708 6503 15714
rect 12434 15708 12486 15714
rect 6503 15665 12434 15699
rect 6451 15650 6503 15656
rect 12434 15650 12486 15656
rect 6727 15631 6779 15637
rect 13131 15631 13183 15637
rect 6779 15588 13131 15622
rect 6727 15573 6779 15579
rect 13131 15573 13183 15579
rect 7003 15554 7055 15560
rect 11092 15554 11144 15560
rect 7055 15511 11092 15545
rect 7003 15496 7055 15502
rect 11092 15496 11144 15502
rect 7279 15477 7331 15483
rect 11789 15477 11841 15483
rect 7331 15434 11789 15468
rect 7279 15419 7331 15425
rect 11789 15419 11841 15425
rect 7555 15400 7607 15406
rect 9750 15400 9802 15406
rect 7607 15357 9750 15391
rect 7555 15342 7607 15348
rect 9750 15342 9802 15348
rect 7831 15323 7883 15329
rect 10447 15323 10499 15329
rect 7883 15280 10447 15314
rect 7831 15265 7883 15271
rect 10447 15265 10499 15271
rect 8107 15246 8159 15252
rect 8482 15246 8534 15252
rect 8159 15203 8482 15237
rect 8107 15188 8159 15194
rect 8482 15188 8534 15194
rect 8383 15169 8435 15175
rect 9105 15169 9157 15175
rect 8435 15126 9105 15160
rect 8383 15111 8435 15117
rect 9105 15111 9157 15117
rect 7140 15092 7192 15098
rect 8659 15092 8711 15098
rect 7192 15049 8659 15083
rect 7140 15034 7192 15040
rect 8659 15034 8711 15040
rect 7689 15015 7741 15021
rect 8935 15015 8987 15021
rect 7741 14972 8935 15006
rect 7689 14957 7741 14963
rect 8935 14957 8987 14963
rect 4382 14938 4434 14944
rect 5724 14938 5776 14944
rect 4434 14895 5510 14929
rect 4382 14880 4434 14886
rect 5079 14861 5131 14867
rect 5131 14818 5433 14852
rect 5079 14803 5131 14809
rect 5399 14698 5433 14818
rect 5476 14775 5510 14895
rect 9211 14938 9263 14944
rect 5776 14895 9211 14929
rect 5724 14880 5776 14886
rect 9211 14880 9263 14886
rect 6347 14861 6399 14867
rect 9487 14861 9539 14867
rect 6399 14818 9487 14852
rect 6347 14803 6399 14809
rect 9487 14803 9539 14809
rect 9763 14784 9815 14790
rect 5476 14741 9763 14775
rect 9763 14726 9815 14732
rect 10039 14707 10091 14713
rect 5399 14664 10039 14698
rect 10039 14649 10091 14655
rect 7729 6940 7781 6946
rect 8163 6940 8215 6946
rect 7781 6897 8163 6931
rect 7729 6882 7781 6888
rect 8163 6882 8215 6888
rect 963 6863 1015 6869
rect 5521 6863 5573 6869
rect 1015 6820 5521 6854
rect 963 6805 1015 6811
rect 5521 6805 5573 6811
rect 8005 6863 8057 6869
rect 8986 6863 9038 6869
rect 8057 6820 8986 6854
rect 8005 6805 8057 6811
rect 8986 6805 9038 6811
rect 1863 6786 1915 6792
rect 5797 6786 5849 6792
rect 1915 6743 5797 6777
rect 1863 6728 1915 6734
rect 5797 6728 5849 6734
rect 8281 6786 8333 6792
rect 10040 6786 10092 6792
rect 8333 6743 10040 6777
rect 8281 6728 8333 6734
rect 10040 6728 10092 6734
rect 2763 6709 2815 6715
rect 6073 6709 6125 6715
rect 2815 6666 6073 6700
rect 2763 6651 2815 6657
rect 6073 6651 6125 6657
rect 8557 6709 8609 6715
rect 10863 6709 10915 6715
rect 8609 6666 10863 6700
rect 8557 6651 8609 6657
rect 10863 6651 10915 6657
rect 3663 6632 3715 6638
rect 6349 6632 6401 6638
rect 3715 6589 6349 6623
rect 3663 6574 3715 6580
rect 6349 6574 6401 6580
rect 8833 6632 8885 6638
rect 11763 6632 11815 6638
rect 8885 6589 11763 6623
rect 8833 6574 8885 6580
rect 11763 6574 11815 6580
rect 4563 6555 4615 6561
rect 6625 6555 6677 6561
rect 4615 6512 6625 6546
rect 4563 6497 4615 6503
rect 6625 6497 6677 6503
rect 9109 6555 9161 6561
rect 12663 6555 12715 6561
rect 9161 6512 12663 6546
rect 9109 6497 9161 6503
rect 12663 6497 12715 6503
rect 5463 6478 5515 6484
rect 6901 6478 6953 6484
rect 5515 6435 6901 6469
rect 5463 6420 5515 6426
rect 6901 6420 6953 6426
rect 9385 6478 9437 6484
rect 13563 6478 13615 6484
rect 9437 6435 13563 6469
rect 9385 6420 9437 6426
rect 13563 6420 13615 6426
rect 6363 6401 6415 6407
rect 7177 6401 7229 6407
rect 6415 6358 7177 6392
rect 6363 6343 6415 6349
rect 7177 6343 7229 6349
rect 9661 6401 9713 6407
rect 14463 6401 14515 6407
rect 9713 6358 14463 6392
rect 9661 6343 9713 6349
rect 14463 6343 14515 6349
rect 7263 6324 7315 6330
rect 7453 6324 7505 6330
rect 7315 6281 7453 6315
rect 7263 6266 7315 6272
rect 7453 6266 7505 6272
rect 9937 6324 9989 6330
rect 15363 6324 15415 6330
rect 9989 6281 15363 6315
rect 9937 6266 9989 6272
rect 15363 6266 15415 6272
rect 963 6038 1015 6044
rect 963 5980 1015 5986
rect 1863 6038 1915 6044
rect 1863 5980 1915 5986
rect 2763 6038 2815 6044
rect 2763 5980 2815 5986
rect 3663 6038 3715 6044
rect 3663 5980 3715 5986
rect 4563 6038 4615 6044
rect 4563 5980 4615 5986
rect 5463 6038 5515 6044
rect 5463 5980 5515 5986
rect 6363 6038 6415 6044
rect 6363 5980 6415 5986
rect 7263 6038 7315 6044
rect 7263 5980 7315 5986
rect 8163 6038 8215 6044
rect 8163 5980 8215 5986
rect 9063 6038 9115 6044
rect 9063 5980 9115 5986
rect 9963 6038 10015 6044
rect 9963 5980 10015 5986
rect 10863 6038 10915 6044
rect 10863 5980 10915 5986
rect 11763 6038 11815 6044
rect 11763 5980 11815 5986
rect 12663 6038 12715 6044
rect 12663 5980 12715 5986
rect 13563 6038 13615 6044
rect 13563 5980 13615 5986
rect 14463 6038 14515 6044
rect 14463 5980 14515 5986
rect 15363 6038 15415 6044
rect 15363 5980 15415 5986
<< via1 >>
rect 4813 20378 4865 20430
rect 7509 20378 7561 20430
rect 10205 20378 10257 20430
rect 12601 20384 12653 20436
rect 12901 20378 12953 20430
rect 5899 15810 5951 15862
rect 13776 15810 13828 15862
rect 6175 15733 6227 15785
rect 14473 15733 14525 15785
rect 6451 15656 6503 15708
rect 12434 15656 12486 15708
rect 6727 15579 6779 15631
rect 13131 15579 13183 15631
rect 7003 15502 7055 15554
rect 11092 15502 11144 15554
rect 7279 15425 7331 15477
rect 11789 15425 11841 15477
rect 7555 15348 7607 15400
rect 9750 15348 9802 15400
rect 7831 15271 7883 15323
rect 10447 15271 10499 15323
rect 8107 15194 8159 15246
rect 8482 15194 8534 15246
rect 8383 15117 8435 15169
rect 9105 15117 9157 15169
rect 7140 15040 7192 15092
rect 8659 15040 8711 15092
rect 7689 14963 7741 15015
rect 8935 14963 8987 15015
rect 4382 14886 4434 14938
rect 5079 14809 5131 14861
rect 5724 14886 5776 14938
rect 9211 14886 9263 14938
rect 6347 14809 6399 14861
rect 9487 14809 9539 14861
rect 9763 14732 9815 14784
rect 10039 14655 10091 14707
rect 7729 6888 7781 6940
rect 8163 6888 8215 6940
rect 963 6811 1015 6863
rect 5521 6811 5573 6863
rect 8005 6811 8057 6863
rect 8986 6811 9038 6863
rect 1863 6734 1915 6786
rect 5797 6734 5849 6786
rect 8281 6734 8333 6786
rect 10040 6734 10092 6786
rect 2763 6657 2815 6709
rect 6073 6657 6125 6709
rect 8557 6657 8609 6709
rect 10863 6657 10915 6709
rect 3663 6580 3715 6632
rect 6349 6580 6401 6632
rect 8833 6580 8885 6632
rect 11763 6580 11815 6632
rect 4563 6503 4615 6555
rect 6625 6503 6677 6555
rect 9109 6503 9161 6555
rect 12663 6503 12715 6555
rect 5463 6426 5515 6478
rect 6901 6426 6953 6478
rect 9385 6426 9437 6478
rect 13563 6426 13615 6478
rect 6363 6349 6415 6401
rect 7177 6349 7229 6401
rect 9661 6349 9713 6401
rect 14463 6349 14515 6401
rect 7263 6272 7315 6324
rect 7453 6272 7505 6324
rect 9937 6272 9989 6324
rect 15363 6272 15415 6324
rect 963 5986 1015 6038
rect 1863 5986 1915 6038
rect 2763 5986 2815 6038
rect 3663 5986 3715 6038
rect 4563 5986 4615 6038
rect 5463 5986 5515 6038
rect 6363 5986 6415 6038
rect 7263 5986 7315 6038
rect 8163 5986 8215 6038
rect 9063 5986 9115 6038
rect 9963 5986 10015 6038
rect 10863 5986 10915 6038
rect 11763 5986 11815 6038
rect 12663 5986 12715 6038
rect 13563 5986 13615 6038
rect 14463 5986 14515 6038
rect 15363 5986 15415 6038
<< metal2 >>
rect 16632 21035 16688 21044
rect 4822 20990 16632 21024
rect 490 19787 499 19977
rect 689 19787 698 19977
rect 564 18655 624 19787
rect 864 19577 924 20467
rect 4822 20436 4856 20990
rect 16632 20970 16688 20979
rect 16506 20953 16562 20962
rect 7518 20908 16506 20942
rect 7518 20436 7552 20908
rect 16506 20888 16562 20897
rect 16884 20871 16940 20880
rect 10214 20826 16884 20860
rect 10214 20436 10248 20826
rect 16884 20806 16940 20815
rect 16380 20789 16436 20798
rect 12610 20744 16380 20778
rect 12610 20442 12644 20744
rect 16380 20724 16436 20733
rect 16758 20707 16814 20716
rect 12910 20662 16758 20696
rect 12601 20436 12653 20442
rect 12910 20436 12944 20662
rect 16758 20642 16814 20651
rect 4813 20430 4865 20436
rect 4813 20372 4865 20378
rect 7509 20430 7561 20436
rect 7509 20372 7561 20378
rect 10205 20430 10257 20436
rect 12601 20378 12653 20384
rect 12901 20430 12953 20436
rect 10205 20372 10257 20378
rect 12901 20372 12953 20378
rect 14672 19577 14732 20467
rect 14898 19787 14907 19977
rect 15097 19787 15106 19977
rect 790 19387 799 19577
rect 989 19387 998 19577
rect 14599 19387 14608 19577
rect 14798 19387 14807 19577
rect 864 18355 924 19387
rect 14672 18355 14732 19387
rect 14972 18655 15032 19787
rect 564 15577 624 16799
rect 488 15387 497 15577
rect 687 15387 696 15577
rect 864 15177 924 17099
rect 790 14987 799 15177
rect 989 14987 998 15177
rect 4391 14938 4425 15982
rect 4769 14987 4778 15177
rect 4968 14987 4977 15177
rect 4376 14886 4382 14938
rect 4434 14886 4440 14938
rect 4823 14686 4923 14987
rect 5088 14861 5122 15982
rect 5273 15387 5282 15577
rect 5472 15387 5481 15577
rect 5073 14809 5079 14861
rect 5131 14809 5137 14861
rect 5327 14686 5427 15387
rect 5733 14938 5767 15982
rect 5893 15810 5899 15862
rect 5951 15810 5957 15862
rect 5718 14886 5724 14938
rect 5776 14886 5782 14938
rect 4823 14586 4995 14686
rect 4895 14384 4995 14586
rect 5045 14586 5427 14686
rect 5045 14384 5145 14586
rect 5908 14572 5942 15810
rect 6169 15733 6175 15785
rect 6227 15733 6233 15785
rect 6430 15776 6464 15982
rect 6356 15742 6464 15776
rect 6184 14572 6218 15733
rect 6356 14861 6390 15742
rect 6445 15656 6451 15708
rect 6503 15656 6509 15708
rect 6341 14809 6347 14861
rect 6399 14809 6405 14861
rect 6460 14572 6494 15656
rect 6721 15579 6727 15631
rect 6779 15579 6785 15631
rect 7075 15622 7109 15982
rect 7075 15588 7183 15622
rect 6736 14572 6770 15579
rect 6997 15502 7003 15554
rect 7055 15502 7061 15554
rect 7012 14572 7046 15502
rect 7149 15092 7183 15588
rect 7273 15425 7279 15477
rect 7331 15425 7337 15477
rect 7134 15040 7140 15092
rect 7192 15040 7198 15092
rect 7288 14572 7322 15425
rect 7549 15348 7555 15400
rect 7607 15348 7613 15400
rect 7772 15391 7806 15982
rect 7698 15357 7806 15391
rect 7564 14572 7598 15348
rect 7698 15015 7732 15357
rect 7825 15271 7831 15323
rect 7883 15271 7889 15323
rect 8417 15314 8451 15982
rect 8417 15280 8525 15314
rect 7683 14963 7689 15015
rect 7741 14963 7747 15015
rect 7840 14572 7874 15271
rect 8491 15246 8525 15280
rect 8101 15194 8107 15246
rect 8159 15194 8165 15246
rect 8476 15194 8482 15246
rect 8534 15194 8540 15246
rect 8116 14572 8150 15194
rect 9114 15169 9148 15982
rect 9759 15400 9793 15982
rect 9744 15348 9750 15400
rect 9802 15348 9808 15400
rect 10164 15387 10173 15577
rect 10363 15387 10372 15577
rect 8377 15117 8383 15169
rect 8435 15117 8441 15169
rect 9099 15117 9105 15169
rect 9157 15117 9163 15169
rect 8392 14572 8426 15117
rect 8653 15040 8659 15092
rect 8711 15040 8717 15092
rect 8668 14572 8702 15040
rect 8929 14963 8935 15015
rect 8987 14963 8993 15015
rect 8944 14572 8978 14963
rect 9205 14886 9211 14938
rect 9263 14886 9269 14938
rect 10218 14886 10318 15387
rect 10456 15323 10490 15982
rect 11101 15554 11135 15982
rect 11086 15502 11092 15554
rect 11144 15502 11150 15554
rect 11798 15477 11832 15982
rect 12443 15708 12477 15982
rect 12428 15656 12434 15708
rect 12486 15656 12492 15708
rect 13140 15631 13174 15982
rect 13785 15862 13819 15982
rect 13770 15810 13776 15862
rect 13828 15810 13834 15862
rect 14482 15785 14516 15982
rect 14467 15733 14473 15785
rect 14525 15733 14531 15785
rect 13125 15579 13131 15631
rect 13183 15579 13189 15631
rect 11783 15425 11789 15477
rect 11841 15425 11847 15477
rect 10441 15271 10447 15323
rect 10499 15271 10505 15323
rect 14672 15177 14732 17099
rect 14972 15577 15032 16799
rect 14897 15387 14906 15577
rect 15096 15387 15105 15577
rect 10565 14987 10574 15177
rect 10764 14987 10773 15177
rect 14599 14987 14608 15177
rect 14798 14987 14807 15177
rect 9220 14572 9254 14886
rect 9481 14809 9487 14861
rect 9539 14809 9545 14861
rect 9496 14572 9530 14809
rect 10218 14786 10567 14886
rect 9757 14732 9763 14784
rect 9815 14732 9821 14784
rect 9772 14572 9806 14732
rect 10033 14655 10039 14707
rect 10091 14655 10097 14707
rect 10048 14572 10082 14655
rect 5888 14516 5897 14572
rect 5953 14516 5962 14572
rect 6164 14516 6173 14572
rect 6229 14516 6238 14572
rect 6440 14516 6449 14572
rect 6505 14516 6514 14572
rect 6716 14516 6725 14572
rect 6781 14516 6790 14572
rect 6992 14516 7001 14572
rect 7057 14516 7066 14572
rect 7268 14516 7277 14572
rect 7333 14516 7342 14572
rect 7544 14516 7553 14572
rect 7609 14516 7618 14572
rect 7820 14516 7829 14572
rect 7885 14516 7894 14572
rect 8096 14516 8105 14572
rect 8161 14516 8170 14572
rect 8372 14516 8381 14572
rect 8437 14516 8446 14572
rect 8648 14516 8657 14572
rect 8713 14516 8722 14572
rect 8924 14516 8933 14572
rect 8989 14516 8998 14572
rect 9200 14516 9209 14572
rect 9265 14516 9274 14572
rect 9476 14516 9485 14572
rect 9541 14516 9550 14572
rect 9752 14516 9761 14572
rect 9817 14516 9826 14572
rect 10028 14516 10037 14572
rect 10093 14516 10102 14572
rect 10467 14384 10567 14786
rect 10617 14384 10717 14987
rect 5895 14237 5955 14246
rect 5895 14010 5955 14181
rect 6171 14237 6231 14246
rect 6171 14010 6231 14181
rect 6447 14237 6507 14246
rect 6447 14010 6507 14181
rect 6723 14237 6783 14246
rect 6723 14010 6783 14181
rect 6999 14237 7059 14246
rect 6999 14010 7059 14181
rect 7275 14237 7335 14246
rect 7275 14010 7335 14181
rect 7551 14237 7611 14246
rect 7551 14010 7611 14181
rect 7827 14237 7887 14246
rect 7827 14010 7887 14181
rect 8103 14237 8163 14246
rect 8103 14010 8163 14181
rect 8379 14237 8439 14246
rect 8379 14010 8439 14181
rect 8655 14237 8715 14246
rect 8655 14010 8715 14181
rect 8931 14237 8991 14246
rect 8931 14010 8991 14181
rect 9207 14237 9267 14246
rect 9207 14010 9267 14181
rect 9483 14237 9543 14246
rect 9483 14010 9543 14181
rect 9759 14237 9819 14246
rect 9759 14010 9819 14181
rect 10035 14237 10095 14246
rect 10035 14010 10095 14181
rect 5517 7393 5577 7562
rect 5517 7328 5577 7337
rect 5793 7393 5853 7562
rect 5793 7328 5853 7337
rect 6069 7393 6129 7562
rect 6069 7328 6129 7337
rect 6345 7393 6405 7562
rect 6345 7328 6405 7337
rect 6621 7393 6681 7562
rect 6621 7328 6681 7337
rect 6897 7393 6957 7562
rect 6897 7328 6957 7337
rect 7173 7393 7233 7562
rect 7173 7328 7233 7337
rect 7449 7393 7509 7562
rect 7449 7328 7509 7337
rect 7725 7393 7785 7562
rect 7725 7328 7785 7337
rect 8001 7393 8061 7562
rect 8001 7328 8061 7337
rect 8277 7393 8337 7562
rect 8277 7328 8337 7337
rect 8553 7393 8613 7562
rect 8553 7328 8613 7337
rect 8829 7393 8889 7562
rect 8829 7328 8889 7337
rect 9105 7393 9165 7562
rect 9105 7328 9165 7337
rect 9381 7393 9441 7562
rect 9381 7328 9441 7337
rect 9657 7393 9717 7562
rect 9657 7328 9717 7337
rect 9933 7393 9993 7562
rect 9933 7328 9993 7337
rect 4840 7088 4995 7188
rect 957 6811 963 6863
rect 1015 6811 1021 6863
rect -4 6405 5 6595
rect 195 6405 204 6595
rect 65 4432 125 6405
rect 972 6038 1006 6811
rect 1857 6734 1863 6786
rect 1915 6734 1921 6786
rect 957 5986 963 6038
rect 1015 5986 1021 6038
rect 1204 6005 1213 6195
rect 1403 6005 1412 6195
rect 1872 6038 1906 6734
rect 2757 6657 2763 6709
rect 2815 6657 2821 6709
rect 2772 6038 2806 6657
rect 3657 6580 3663 6632
rect 3715 6580 3721 6632
rect 3672 6038 3706 6580
rect 4557 6503 4563 6555
rect 4615 6503 4621 6555
rect 4572 6038 4606 6503
rect 4840 6195 4940 7088
rect 5045 6595 5145 7188
rect 5510 7004 5519 7060
rect 5575 7004 5584 7060
rect 5786 7004 5795 7060
rect 5851 7004 5860 7060
rect 6062 7004 6071 7060
rect 6127 7004 6136 7060
rect 6338 7004 6347 7060
rect 6403 7004 6412 7060
rect 6614 7004 6623 7060
rect 6679 7004 6688 7060
rect 6890 7004 6899 7060
rect 6955 7004 6964 7060
rect 7166 7004 7175 7060
rect 7231 7004 7240 7060
rect 7442 7004 7451 7060
rect 7507 7004 7516 7060
rect 7718 7004 7727 7060
rect 7783 7004 7792 7060
rect 7994 7004 8003 7060
rect 8059 7004 8068 7060
rect 8270 7004 8279 7060
rect 8335 7004 8344 7060
rect 8546 7004 8555 7060
rect 8611 7004 8620 7060
rect 8822 7004 8831 7060
rect 8887 7004 8896 7060
rect 9098 7004 9107 7060
rect 9163 7004 9172 7060
rect 9374 7004 9383 7060
rect 9439 7004 9448 7060
rect 9650 7004 9659 7060
rect 9715 7004 9724 7060
rect 9926 7004 9935 7060
rect 9991 7004 10000 7060
rect 5530 6863 5564 7004
rect 5515 6811 5521 6863
rect 5573 6811 5579 6863
rect 5806 6786 5840 7004
rect 5791 6734 5797 6786
rect 5849 6734 5855 6786
rect 6082 6709 6116 7004
rect 6067 6657 6073 6709
rect 6125 6657 6131 6709
rect 6358 6632 6392 7004
rect 4989 6405 4998 6595
rect 5188 6405 5197 6595
rect 6343 6580 6349 6632
rect 6401 6580 6407 6632
rect 6634 6555 6668 7004
rect 6619 6503 6625 6555
rect 6677 6503 6683 6555
rect 6910 6478 6944 7004
rect 5457 6426 5463 6478
rect 5515 6426 5521 6478
rect 6895 6426 6901 6478
rect 6953 6426 6959 6478
rect 1278 5815 1338 6005
rect 1857 5986 1863 6038
rect 1915 5986 1921 6038
rect 2757 5986 2763 6038
rect 2815 5986 2821 6038
rect 3657 5986 3663 6038
rect 3715 5986 3721 6038
rect 4557 5986 4563 6038
rect 4615 5986 4621 6038
rect 4786 6005 4795 6195
rect 4985 6005 4994 6195
rect 5472 6038 5506 6426
rect 7186 6401 7220 7004
rect 6357 6349 6363 6401
rect 6415 6349 6421 6401
rect 7171 6349 7177 6401
rect 7229 6349 7235 6401
rect 6372 6038 6406 6349
rect 7462 6324 7496 7004
rect 7738 6940 7772 7004
rect 7723 6888 7729 6940
rect 7781 6888 7787 6940
rect 8014 6863 8048 7004
rect 8157 6888 8163 6940
rect 8215 6888 8221 6940
rect 7999 6811 8005 6863
rect 8057 6811 8063 6863
rect 7257 6272 7263 6324
rect 7315 6272 7321 6324
rect 7447 6272 7453 6324
rect 7505 6272 7511 6324
rect 7272 6038 7306 6272
rect 8172 6038 8206 6888
rect 8290 6786 8324 7004
rect 8275 6734 8281 6786
rect 8333 6734 8339 6786
rect 8566 6709 8600 7004
rect 8551 6657 8557 6709
rect 8609 6657 8615 6709
rect 8842 6632 8876 7004
rect 8980 6811 8986 6863
rect 9038 6811 9044 6863
rect 8827 6580 8833 6632
rect 8885 6580 8891 6632
rect 8995 6190 9029 6811
rect 9118 6555 9152 7004
rect 9103 6503 9109 6555
rect 9161 6503 9167 6555
rect 9394 6478 9428 7004
rect 9379 6426 9385 6478
rect 9437 6426 9443 6478
rect 9670 6401 9704 7004
rect 9655 6349 9661 6401
rect 9713 6349 9719 6401
rect 9946 6324 9980 7004
rect 10467 6988 10567 7188
rect 10366 6888 10567 6988
rect 10034 6734 10040 6786
rect 10092 6734 10098 6786
rect 9931 6272 9937 6324
rect 9989 6272 9995 6324
rect 10049 6190 10083 6734
rect 10366 6595 10466 6888
rect 10312 6405 10321 6595
rect 10511 6405 10520 6595
rect 10617 6195 10717 7188
rect 10857 6657 10863 6709
rect 10915 6657 10921 6709
rect 8995 6156 9106 6190
rect 9072 6038 9106 6156
rect 9972 6156 10083 6190
rect 9972 6038 10006 6156
rect 5457 5986 5463 6038
rect 5515 5986 5521 6038
rect 6357 5986 6363 6038
rect 6415 5986 6421 6038
rect 7257 5986 7263 6038
rect 7315 5986 7321 6038
rect 8157 5986 8163 6038
rect 8215 5986 8221 6038
rect 9057 5986 9063 6038
rect 9115 5986 9121 6038
rect 9957 5986 9963 6038
rect 10015 5986 10021 6038
rect 10564 6005 10573 6195
rect 10763 6005 10772 6195
rect 10872 6038 10906 6657
rect 11757 6580 11763 6632
rect 11815 6580 11821 6632
rect 11772 6038 11806 6580
rect 12657 6503 12663 6555
rect 12715 6503 12721 6555
rect 12672 6038 12706 6503
rect 13557 6426 13563 6478
rect 13615 6426 13621 6478
rect 13572 6038 13606 6426
rect 15392 6405 15401 6595
rect 15591 6405 15600 6595
rect 14457 6349 14463 6401
rect 14515 6349 14521 6401
rect 14472 6038 14506 6349
rect 15357 6272 15363 6324
rect 15415 6272 15421 6324
rect 10857 5986 10863 6038
rect 10915 5986 10921 6038
rect 11757 5986 11763 6038
rect 11815 5986 11821 6038
rect 12657 5986 12663 6038
rect 12715 5986 12721 6038
rect 13557 5986 13563 6038
rect 13615 5986 13621 6038
rect 14457 5986 14463 6038
rect 14515 5986 14521 6038
rect 14748 6005 14757 6195
rect 14947 6005 14956 6195
rect 15372 6038 15406 6272
rect 14823 5826 14883 6005
rect 15357 5986 15363 6038
rect 15415 5986 15421 6038
rect 1056 5755 1338 5815
rect 14570 5766 14883 5826
rect 1056 5382 1116 5755
rect 899 5322 1116 5382
rect 14570 5382 14630 5766
rect 14570 5322 14883 5382
rect 899 3072 959 5322
rect 14823 4895 14883 5322
rect 14823 4835 15067 4895
rect 15007 4518 15067 4835
rect 15471 4432 15531 6405
rect 599 595 659 1516
rect 523 405 532 595
rect 722 405 731 595
rect 899 195 959 1816
rect 826 5 835 195
rect 1025 5 1034 195
rect 9864 -342 9898 434
rect 11206 -260 11240 438
rect 12548 -178 12582 434
rect 13890 -96 13924 434
rect 15007 195 15067 1816
rect 15307 595 15367 1516
rect 15234 405 15243 595
rect 15433 405 15442 595
rect 14932 5 14941 195
rect 15131 5 15140 195
rect 16128 -85 16184 -76
rect 13890 -130 16128 -96
rect 16128 -150 16184 -141
rect 16002 -167 16058 -158
rect 12548 -212 16002 -178
rect 16002 -232 16058 -223
rect 16380 -249 16436 -240
rect 11206 -294 16380 -260
rect 16380 -314 16436 -305
rect 16254 -331 16310 -322
rect 9864 -376 16254 -342
rect 16254 -396 16310 -387
<< via2 >>
rect 499 19787 689 19977
rect 16632 20979 16688 21035
rect 16506 20897 16562 20953
rect 16884 20815 16940 20871
rect 16380 20733 16436 20789
rect 16758 20651 16814 20707
rect 14907 19787 15097 19977
rect 799 19387 989 19577
rect 14608 19387 14798 19577
rect 497 15387 687 15577
rect 799 14987 989 15177
rect 4778 14987 4968 15177
rect 5282 15387 5472 15577
rect 10173 15387 10363 15577
rect 14906 15387 15096 15577
rect 10574 14987 10764 15177
rect 14608 14987 14798 15177
rect 5897 14516 5953 14572
rect 6173 14516 6229 14572
rect 6449 14516 6505 14572
rect 6725 14516 6781 14572
rect 7001 14516 7057 14572
rect 7277 14516 7333 14572
rect 7553 14516 7609 14572
rect 7829 14516 7885 14572
rect 8105 14516 8161 14572
rect 8381 14516 8437 14572
rect 8657 14516 8713 14572
rect 8933 14516 8989 14572
rect 9209 14516 9265 14572
rect 9485 14516 9541 14572
rect 9761 14516 9817 14572
rect 10037 14516 10093 14572
rect 5895 14181 5955 14237
rect 6171 14181 6231 14237
rect 6447 14181 6507 14237
rect 6723 14181 6783 14237
rect 6999 14181 7059 14237
rect 7275 14181 7335 14237
rect 7551 14181 7611 14237
rect 7827 14181 7887 14237
rect 8103 14181 8163 14237
rect 8379 14181 8439 14237
rect 8655 14181 8715 14237
rect 8931 14181 8991 14237
rect 9207 14181 9267 14237
rect 9483 14181 9543 14237
rect 9759 14181 9819 14237
rect 10035 14181 10095 14237
rect 5517 7337 5577 7393
rect 5793 7337 5853 7393
rect 6069 7337 6129 7393
rect 6345 7337 6405 7393
rect 6621 7337 6681 7393
rect 6897 7337 6957 7393
rect 7173 7337 7233 7393
rect 7449 7337 7509 7393
rect 7725 7337 7785 7393
rect 8001 7337 8061 7393
rect 8277 7337 8337 7393
rect 8553 7337 8613 7393
rect 8829 7337 8889 7393
rect 9105 7337 9165 7393
rect 9381 7337 9441 7393
rect 9657 7337 9717 7393
rect 9933 7337 9993 7393
rect 5 6405 195 6595
rect 1213 6005 1403 6195
rect 5519 7004 5575 7060
rect 5795 7004 5851 7060
rect 6071 7004 6127 7060
rect 6347 7004 6403 7060
rect 6623 7004 6679 7060
rect 6899 7004 6955 7060
rect 7175 7004 7231 7060
rect 7451 7004 7507 7060
rect 7727 7004 7783 7060
rect 8003 7004 8059 7060
rect 8279 7004 8335 7060
rect 8555 7004 8611 7060
rect 8831 7004 8887 7060
rect 9107 7004 9163 7060
rect 9383 7004 9439 7060
rect 9659 7004 9715 7060
rect 9935 7004 9991 7060
rect 4998 6405 5188 6595
rect 4795 6005 4985 6195
rect 10321 6405 10511 6595
rect 10573 6005 10763 6195
rect 15401 6405 15591 6595
rect 14757 6005 14947 6195
rect 532 405 722 595
rect 835 5 1025 195
rect 15243 405 15433 595
rect 14941 5 15131 195
rect 16128 -141 16184 -85
rect 16002 -223 16058 -167
rect 16380 -305 16436 -249
rect 16254 -387 16310 -331
<< metal3 >>
rect 0 19977 15596 19982
rect 0 19787 499 19977
rect 689 19787 14907 19977
rect 15097 19787 15596 19977
rect 0 19782 15596 19787
rect 0 19577 15596 19582
rect 0 19387 799 19577
rect 989 19387 14608 19577
rect 14798 19387 15596 19577
rect 0 19382 15596 19387
rect 0 15577 15596 15582
rect 0 15387 497 15577
rect 687 15387 5282 15577
rect 5472 15387 10173 15577
rect 10363 15387 14906 15577
rect 15096 15387 15596 15577
rect 0 15382 15596 15387
rect 0 15177 15596 15182
rect 0 14987 799 15177
rect 989 14987 4778 15177
rect 4968 14987 10574 15177
rect 10764 14987 14608 15177
rect 14798 14987 15596 15177
rect 0 14982 15596 14987
rect 5892 14572 5958 14577
rect 5892 14516 5897 14572
rect 5953 14516 5958 14572
rect 5892 14511 5958 14516
rect 6168 14572 6234 14577
rect 6168 14516 6173 14572
rect 6229 14516 6234 14572
rect 6168 14511 6234 14516
rect 6444 14572 6510 14577
rect 6444 14516 6449 14572
rect 6505 14516 6510 14572
rect 6444 14511 6510 14516
rect 6720 14572 6786 14577
rect 6720 14516 6725 14572
rect 6781 14516 6786 14572
rect 6720 14511 6786 14516
rect 6996 14572 7062 14577
rect 6996 14516 7001 14572
rect 7057 14516 7062 14572
rect 6996 14511 7062 14516
rect 7272 14572 7338 14577
rect 7272 14516 7277 14572
rect 7333 14516 7338 14572
rect 7272 14511 7338 14516
rect 7548 14572 7614 14577
rect 7548 14516 7553 14572
rect 7609 14516 7614 14572
rect 7548 14511 7614 14516
rect 7824 14572 7890 14577
rect 7824 14516 7829 14572
rect 7885 14516 7890 14572
rect 7824 14511 7890 14516
rect 8100 14572 8166 14577
rect 8100 14516 8105 14572
rect 8161 14516 8166 14572
rect 8100 14511 8166 14516
rect 8376 14572 8442 14577
rect 8376 14516 8381 14572
rect 8437 14516 8442 14572
rect 8376 14511 8442 14516
rect 8652 14572 8718 14577
rect 8652 14516 8657 14572
rect 8713 14516 8718 14572
rect 8652 14511 8718 14516
rect 8928 14572 8994 14577
rect 8928 14516 8933 14572
rect 8989 14516 8994 14572
rect 8928 14511 8994 14516
rect 9204 14572 9270 14577
rect 9204 14516 9209 14572
rect 9265 14516 9270 14572
rect 9204 14511 9270 14516
rect 9480 14572 9546 14577
rect 9480 14516 9485 14572
rect 9541 14516 9546 14572
rect 9480 14511 9546 14516
rect 9756 14572 9822 14577
rect 9756 14516 9761 14572
rect 9817 14516 9822 14572
rect 9756 14511 9822 14516
rect 10032 14572 10098 14577
rect 10032 14516 10037 14572
rect 10093 14516 10098 14572
rect 10032 14511 10098 14516
rect 5895 14242 5955 14511
rect 6171 14242 6231 14511
rect 6447 14242 6507 14511
rect 6723 14242 6783 14511
rect 6999 14242 7059 14511
rect 7275 14242 7335 14511
rect 7551 14242 7611 14511
rect 7827 14242 7887 14511
rect 8103 14242 8163 14511
rect 8379 14242 8439 14511
rect 8655 14242 8715 14511
rect 8931 14242 8991 14511
rect 9207 14242 9267 14511
rect 9483 14242 9543 14511
rect 9759 14242 9819 14511
rect 10035 14242 10095 14511
rect 5890 14237 5960 14242
rect 5890 14181 5895 14237
rect 5955 14181 5960 14237
rect 5890 14176 5960 14181
rect 6166 14237 6236 14242
rect 6166 14181 6171 14237
rect 6231 14181 6236 14237
rect 6166 14176 6236 14181
rect 6442 14237 6512 14242
rect 6442 14181 6447 14237
rect 6507 14181 6512 14237
rect 6442 14176 6512 14181
rect 6718 14237 6788 14242
rect 6718 14181 6723 14237
rect 6783 14181 6788 14237
rect 6718 14176 6788 14181
rect 6994 14237 7064 14242
rect 6994 14181 6999 14237
rect 7059 14181 7064 14237
rect 6994 14176 7064 14181
rect 7270 14237 7340 14242
rect 7270 14181 7275 14237
rect 7335 14181 7340 14237
rect 7270 14176 7340 14181
rect 7546 14237 7616 14242
rect 7546 14181 7551 14237
rect 7611 14181 7616 14237
rect 7546 14176 7616 14181
rect 7822 14237 7892 14242
rect 7822 14181 7827 14237
rect 7887 14181 7892 14237
rect 7822 14176 7892 14181
rect 8098 14237 8168 14242
rect 8098 14181 8103 14237
rect 8163 14181 8168 14237
rect 8098 14176 8168 14181
rect 8374 14237 8444 14242
rect 8374 14181 8379 14237
rect 8439 14181 8444 14237
rect 8374 14176 8444 14181
rect 8650 14237 8720 14242
rect 8650 14181 8655 14237
rect 8715 14181 8720 14237
rect 8650 14176 8720 14181
rect 8926 14237 8996 14242
rect 8926 14181 8931 14237
rect 8991 14181 8996 14237
rect 8926 14176 8996 14181
rect 9202 14237 9272 14242
rect 9202 14181 9207 14237
rect 9267 14181 9272 14237
rect 9202 14176 9272 14181
rect 9478 14237 9548 14242
rect 9478 14181 9483 14237
rect 9543 14181 9548 14237
rect 9478 14176 9548 14181
rect 9754 14237 9824 14242
rect 9754 14181 9759 14237
rect 9819 14181 9824 14237
rect 9754 14176 9824 14181
rect 10030 14237 10100 14242
rect 10030 14181 10035 14237
rect 10095 14181 10100 14237
rect 10030 14176 10100 14181
rect 5856 13799 10134 13937
rect 5512 7393 5582 7398
rect 5512 7337 5517 7393
rect 5577 7337 5582 7393
rect 5512 7332 5582 7337
rect 5788 7393 5858 7398
rect 5788 7337 5793 7393
rect 5853 7337 5858 7393
rect 5788 7332 5858 7337
rect 6064 7393 6134 7398
rect 6064 7337 6069 7393
rect 6129 7337 6134 7393
rect 6064 7332 6134 7337
rect 6340 7393 6410 7398
rect 6340 7337 6345 7393
rect 6405 7337 6410 7393
rect 6340 7332 6410 7337
rect 6616 7393 6686 7398
rect 6616 7337 6621 7393
rect 6681 7337 6686 7393
rect 6616 7332 6686 7337
rect 6892 7393 6962 7398
rect 6892 7337 6897 7393
rect 6957 7337 6962 7393
rect 6892 7332 6962 7337
rect 7168 7393 7238 7398
rect 7168 7337 7173 7393
rect 7233 7337 7238 7393
rect 7168 7332 7238 7337
rect 7444 7393 7514 7398
rect 7444 7337 7449 7393
rect 7509 7337 7514 7393
rect 7444 7332 7514 7337
rect 7720 7393 7790 7398
rect 7720 7337 7725 7393
rect 7785 7337 7790 7393
rect 7720 7332 7790 7337
rect 7996 7393 8066 7398
rect 7996 7337 8001 7393
rect 8061 7337 8066 7393
rect 7996 7332 8066 7337
rect 8272 7393 8342 7398
rect 8272 7337 8277 7393
rect 8337 7337 8342 7393
rect 8272 7332 8342 7337
rect 8548 7393 8618 7398
rect 8548 7337 8553 7393
rect 8613 7337 8618 7393
rect 8548 7332 8618 7337
rect 8824 7393 8894 7398
rect 8824 7337 8829 7393
rect 8889 7337 8894 7393
rect 8824 7332 8894 7337
rect 9100 7393 9170 7398
rect 9100 7337 9105 7393
rect 9165 7337 9170 7393
rect 9100 7332 9170 7337
rect 9376 7393 9446 7398
rect 9376 7337 9381 7393
rect 9441 7337 9446 7393
rect 9376 7332 9446 7337
rect 9652 7393 9722 7398
rect 9652 7337 9657 7393
rect 9717 7337 9722 7393
rect 9652 7332 9722 7337
rect 9928 7393 9998 7398
rect 9928 7337 9933 7393
rect 9993 7337 9998 7393
rect 9928 7332 9998 7337
rect 5517 7065 5577 7332
rect 5793 7065 5853 7332
rect 6069 7065 6129 7332
rect 6345 7065 6405 7332
rect 6621 7065 6681 7332
rect 6897 7065 6957 7332
rect 7173 7065 7233 7332
rect 7449 7065 7509 7332
rect 7725 7065 7785 7332
rect 8001 7065 8061 7332
rect 8277 7065 8337 7332
rect 8553 7065 8613 7332
rect 8829 7065 8889 7332
rect 9105 7065 9165 7332
rect 9381 7065 9441 7332
rect 9657 7065 9717 7332
rect 9933 7065 9993 7332
rect 5514 7060 5580 7065
rect 5514 7004 5519 7060
rect 5575 7004 5580 7060
rect 5514 6999 5580 7004
rect 5790 7060 5856 7065
rect 5790 7004 5795 7060
rect 5851 7004 5856 7060
rect 5790 6999 5856 7004
rect 6066 7060 6132 7065
rect 6066 7004 6071 7060
rect 6127 7004 6132 7060
rect 6066 6999 6132 7004
rect 6342 7060 6408 7065
rect 6342 7004 6347 7060
rect 6403 7004 6408 7060
rect 6342 6999 6408 7004
rect 6618 7060 6684 7065
rect 6618 7004 6623 7060
rect 6679 7004 6684 7060
rect 6618 6999 6684 7004
rect 6894 7060 6960 7065
rect 6894 7004 6899 7060
rect 6955 7004 6960 7060
rect 6894 6999 6960 7004
rect 7170 7060 7236 7065
rect 7170 7004 7175 7060
rect 7231 7004 7236 7060
rect 7170 6999 7236 7004
rect 7446 7060 7512 7065
rect 7446 7004 7451 7060
rect 7507 7004 7512 7060
rect 7446 6999 7512 7004
rect 7722 7060 7788 7065
rect 7722 7004 7727 7060
rect 7783 7004 7788 7060
rect 7722 6999 7788 7004
rect 7998 7060 8064 7065
rect 7998 7004 8003 7060
rect 8059 7004 8064 7060
rect 7998 6999 8064 7004
rect 8274 7060 8340 7065
rect 8274 7004 8279 7060
rect 8335 7004 8340 7060
rect 8274 6999 8340 7004
rect 8550 7060 8616 7065
rect 8550 7004 8555 7060
rect 8611 7004 8616 7060
rect 8550 6999 8616 7004
rect 8826 7060 8892 7065
rect 8826 7004 8831 7060
rect 8887 7004 8892 7060
rect 8826 6999 8892 7004
rect 9102 7060 9168 7065
rect 9102 7004 9107 7060
rect 9163 7004 9168 7060
rect 9102 6999 9168 7004
rect 9378 7060 9444 7065
rect 9378 7004 9383 7060
rect 9439 7004 9444 7060
rect 9378 6999 9444 7004
rect 9654 7060 9720 7065
rect 9654 7004 9659 7060
rect 9715 7004 9720 7060
rect 9654 6999 9720 7004
rect 9930 7060 9996 7065
rect 9930 7004 9935 7060
rect 9991 7004 9996 7060
rect 9930 6999 9996 7004
rect 0 6595 15596 6600
rect 0 6405 5 6595
rect 195 6405 4998 6595
rect 5188 6405 10321 6595
rect 10511 6405 15401 6595
rect 15591 6405 15596 6595
rect 0 6400 15596 6405
rect 0 6195 15596 6200
rect 0 6005 1213 6195
rect 1403 6005 4795 6195
rect 4985 6005 10573 6195
rect 10763 6005 14757 6195
rect 14947 6005 15596 6195
rect 0 6000 15596 6005
rect 0 595 15596 600
rect 0 405 532 595
rect 722 405 15243 595
rect 15433 405 15596 595
rect 0 400 15596 405
rect 0 195 15596 200
rect 0 5 835 195
rect 1025 5 14941 195
rect 15131 5 15596 195
rect 0 0 15596 5
rect 16000 -162 16060 21435
rect 16126 -80 16186 21435
rect 16123 -85 16189 -80
rect 16123 -141 16128 -85
rect 16184 -141 16189 -85
rect 16123 -146 16189 -141
rect 15997 -167 16063 -162
rect 15997 -223 16002 -167
rect 16058 -223 16063 -167
rect 15997 -228 16063 -223
rect 16252 -326 16312 21435
rect 16378 20794 16438 21435
rect 16504 20958 16564 21435
rect 16630 21040 16690 21435
rect 16627 21035 16693 21040
rect 16627 20979 16632 21035
rect 16688 20979 16693 21035
rect 16627 20974 16693 20979
rect 16501 20953 16567 20958
rect 16501 20897 16506 20953
rect 16562 20897 16567 20953
rect 16501 20892 16567 20897
rect 16375 20789 16441 20794
rect 16375 20733 16380 20789
rect 16436 20733 16441 20789
rect 16375 20728 16441 20733
rect 16378 -244 16438 20728
rect 16504 0 16564 20892
rect 16756 20712 16816 21435
rect 16882 20876 16942 21435
rect 16879 20871 16945 20876
rect 16879 20815 16884 20871
rect 16940 20815 16945 20871
rect 16879 20810 16945 20815
rect 16753 20707 16819 20712
rect 16753 20651 16758 20707
rect 16814 20651 16819 20707
rect 16753 20646 16819 20651
rect 16375 -249 16441 -244
rect 16375 -305 16380 -249
rect 16436 -305 16441 -249
rect 16375 -310 16441 -305
rect 16249 -331 16315 -326
rect 16249 -387 16254 -331
rect 16310 -387 16315 -331
rect 16249 -392 16315 -387
use dac_main  dac_main_0
timestamp 1748337984
transform 1 0 4895 0 1 7088
box 0 0 5822 7396
use lsb_decoder  lsb_decoder_0
timestamp 1748337480
transform 1 0 1128 0 1 15870
box -571 0 13911 4692
use msb_decoder  msb_decoder_0
timestamp 1748318706
transform 1 0 0 0 1 400
box 0 0 15596 5868
<< labels >>
flabel metal3 0 0 15596 200 0 FreeSans 256 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 0 400 15596 600 0 FreeSans 256 0 0 0 VDD
port 2 nsew power bidirectional
flabel metal3 5856 13799 10134 13937 0 FreeSans 256 0 0 0 VOUT
port 3 nsew signal bidirectional
flabel metal3 16882 21135 16942 21435 0 FreeSans 256 0 0 0 IN[0]
port 4 nsew signal input
flabel metal3 16756 21135 16816 21435 0 FreeSans 256 0 0 0 IN[1]
port 5 nsew signal input
flabel metal3 16630 21135 16690 21435 0 FreeSans 256 0 0 0 IN[2]
port 6 nsew signal input
flabel metal3 16504 21135 16564 21435 0 FreeSans 256 0 0 0 IN[3]
port 7 nsew signal input
flabel metal3 16378 21135 16438 21435 0 FreeSans 256 0 0 0 IN[4]
port 8 nsew signal input
flabel metal3 16252 21135 16312 21435 0 FreeSans 256 0 0 0 IN[5]
port 9 nsew signal input
flabel metal3 16126 21135 16186 21435 0 FreeSans 256 0 0 0 IN[6]
port 10 nsew signal input
flabel metal3 16000 21135 16060 21435 0 FreeSans 256 0 0 0 IN[7]
port 11 nsew signal input
<< end >>
