magic
tech sky130A
magscale 1 2
timestamp 1748318706
<< viali >>
rect 78 5356 112 5694
rect 15484 5356 15518 5694
rect 58 4720 92 4988
rect 15514 4720 15548 4988
<< metal1 >>
rect 63 5703 127 5709
rect 63 5347 69 5703
rect 121 5347 127 5703
rect 15469 5703 15533 5709
rect 63 5341 127 5347
rect 45 4988 105 5001
rect 45 4720 58 4988
rect 92 4720 105 4988
rect 972 4785 1006 5629
rect 1872 4785 1906 5629
rect 2772 4785 2806 5629
rect 3672 4785 3706 5629
rect 4572 4785 4606 5629
rect 5472 4785 5506 5629
rect 6372 4785 6406 5629
rect 7272 4785 7306 5629
rect 8172 4785 8206 5629
rect 9072 4785 9106 5629
rect 9972 4785 10006 5629
rect 10872 4785 10906 5629
rect 11772 4785 11806 5629
rect 12672 4785 12706 5629
rect 13572 4785 13606 5629
rect 14472 4785 14506 5629
rect 15372 4785 15406 5629
rect 15469 5347 15475 5703
rect 15527 5347 15533 5703
rect 15469 5341 15533 5347
rect 15501 4988 15561 5001
rect 45 4392 105 4720
rect 272 4760 324 4766
rect 272 4702 324 4708
rect 572 4760 624 4766
rect 572 4702 624 4708
rect 1172 4760 1224 4766
rect 1172 4702 1224 4708
rect 1472 4760 1524 4766
rect 1472 4702 1524 4708
rect 2072 4760 2124 4766
rect 2072 4702 2124 4708
rect 2372 4760 2424 4766
rect 2372 4702 2424 4708
rect 2972 4760 3024 4766
rect 2972 4702 3024 4708
rect 3272 4760 3324 4766
rect 3272 4702 3324 4708
rect 3872 4760 3924 4766
rect 3872 4702 3924 4708
rect 4172 4760 4224 4766
rect 4172 4702 4224 4708
rect 4772 4760 4824 4766
rect 4772 4702 4824 4708
rect 5072 4760 5124 4766
rect 5072 4702 5124 4708
rect 5672 4760 5724 4766
rect 5672 4702 5724 4708
rect 5972 4760 6024 4766
rect 5972 4702 6024 4708
rect 6572 4760 6624 4766
rect 6572 4702 6624 4708
rect 6872 4760 6924 4766
rect 6872 4702 6924 4708
rect 7472 4760 7524 4766
rect 7472 4702 7524 4708
rect 7772 4760 7824 4766
rect 7772 4702 7824 4708
rect 8372 4760 8424 4766
rect 8372 4702 8424 4708
rect 8672 4760 8724 4766
rect 8672 4702 8724 4708
rect 9272 4760 9324 4766
rect 9272 4702 9324 4708
rect 9572 4760 9624 4766
rect 9572 4702 9624 4708
rect 10172 4760 10224 4766
rect 10172 4702 10224 4708
rect 10472 4760 10524 4766
rect 10472 4702 10524 4708
rect 11072 4760 11124 4766
rect 11072 4702 11124 4708
rect 11372 4760 11424 4766
rect 11372 4702 11424 4708
rect 11972 4760 12024 4766
rect 11972 4702 12024 4708
rect 12272 4760 12324 4766
rect 12272 4702 12324 4708
rect 12872 4760 12924 4766
rect 12872 4702 12924 4708
rect 13172 4760 13224 4766
rect 13172 4702 13224 4708
rect 13772 4760 13824 4766
rect 13772 4702 13824 4708
rect 14072 4760 14124 4766
rect 14072 4702 14124 4708
rect 14672 4760 14724 4766
rect 14672 4702 14724 4708
rect 14972 4760 15024 4766
rect 14972 4702 15024 4708
rect 15501 4720 15514 4988
rect 15548 4720 15561 4988
rect 272 4667 324 4673
rect 272 4609 324 4615
rect 14972 4667 15024 4673
rect 14972 4609 15024 4615
rect 572 4542 624 4548
rect 1172 4542 1224 4548
rect 624 4499 1172 4533
rect 572 4484 624 4490
rect 10600 4542 10652 4548
rect 1224 4499 10600 4533
rect 1172 4484 1224 4490
rect 10600 4484 10652 4490
rect 1472 4465 1524 4471
rect 2072 4465 2124 4471
rect 1524 4422 2072 4456
rect 1472 4407 1524 4413
rect 11197 4465 11249 4471
rect 2124 4422 11197 4456
rect 2072 4407 2124 4413
rect 11197 4407 11249 4413
rect 899 4392 959 4398
rect 45 4332 899 4392
rect 899 4326 959 4332
rect 2372 4388 2424 4394
rect 2972 4388 3024 4394
rect 2424 4345 2972 4379
rect 2372 4330 2424 4336
rect 9158 4388 9210 4394
rect 3024 4345 9158 4379
rect 2972 4330 3024 4336
rect 9158 4330 9210 4336
rect 15007 4392 15067 4398
rect 15501 4392 15561 4720
rect 15067 4332 15561 4392
rect 15007 4326 15067 4332
rect 3272 4311 3324 4317
rect 3872 4311 3924 4317
rect 3324 4268 3872 4302
rect 3272 4253 3324 4259
rect 9855 4311 9907 4317
rect 3924 4268 9855 4302
rect 3872 4253 3924 4259
rect 9855 4253 9907 4259
rect 4172 4234 4224 4240
rect 4772 4234 4824 4240
rect 4224 4191 4772 4225
rect 4172 4176 4224 4182
rect 7916 4234 7968 4240
rect 4824 4191 7916 4225
rect 4772 4176 4824 4182
rect 7916 4176 7968 4182
rect 5072 4157 5124 4163
rect 5672 4157 5724 4163
rect 5124 4114 5672 4148
rect 5072 4099 5124 4105
rect 8513 4157 8565 4163
rect 5724 4114 8513 4148
rect 5672 4099 5724 4105
rect 8513 4099 8565 4105
rect 5972 4080 6024 4086
rect 6474 4080 6526 4086
rect 6024 4037 6474 4071
rect 5972 4022 6024 4028
rect 6572 4080 6624 4086
rect 6526 4037 6572 4071
rect 6474 4022 6526 4028
rect 6572 4022 6624 4028
rect 6872 4003 6924 4009
rect 7171 4003 7223 4009
rect 6924 3960 7171 3994
rect 6872 3945 6924 3951
rect 7472 4003 7524 4009
rect 7223 3960 7472 3994
rect 7171 3945 7223 3951
rect 7472 3945 7524 3951
rect 5132 3926 5184 3932
rect 7772 3926 7824 3932
rect 5184 3883 7772 3917
rect 5132 3868 5184 3874
rect 8372 3926 8424 3932
rect 7824 3883 8372 3917
rect 7772 3868 7824 3874
rect 8372 3868 8424 3874
rect 5829 3849 5881 3855
rect 8672 3849 8724 3855
rect 5881 3806 8672 3840
rect 5829 3791 5881 3797
rect 9272 3849 9324 3855
rect 8724 3806 9272 3840
rect 8672 3791 8724 3797
rect 9272 3791 9324 3797
rect 3790 3772 3842 3778
rect 9572 3772 9624 3778
rect 3842 3729 9572 3763
rect 3790 3714 3842 3720
rect 10172 3772 10224 3778
rect 9624 3729 10172 3763
rect 9572 3714 9624 3720
rect 10172 3714 10224 3720
rect 4487 3695 4539 3701
rect 10472 3695 10524 3701
rect 4539 3652 10472 3686
rect 4487 3637 4539 3643
rect 11072 3695 11124 3701
rect 10524 3652 11072 3686
rect 10472 3637 10524 3643
rect 11072 3637 11124 3643
rect 2448 3618 2500 3624
rect 11372 3618 11424 3624
rect 2500 3575 11372 3609
rect 2448 3560 2500 3566
rect 11972 3618 12024 3624
rect 11424 3575 11972 3609
rect 11372 3560 11424 3566
rect 11972 3560 12024 3566
rect 3145 3541 3197 3547
rect 12272 3541 12324 3547
rect 3197 3498 12272 3532
rect 3145 3483 3197 3489
rect 12872 3541 12924 3547
rect 12324 3498 12872 3532
rect 12272 3483 12324 3489
rect 12872 3483 12924 3489
rect 1106 3464 1158 3470
rect 13172 3464 13224 3470
rect 1158 3421 13172 3455
rect 1106 3406 1158 3412
rect 13772 3464 13824 3470
rect 13224 3421 13772 3455
rect 13172 3406 13224 3412
rect 13772 3406 13824 3412
rect 1803 3387 1855 3393
rect 14072 3387 14124 3393
rect 1855 3344 14072 3378
rect 1803 3329 1855 3335
rect 14672 3387 14724 3393
rect 14124 3344 14672 3378
rect 14072 3329 14124 3335
rect 14672 3329 14724 3335
<< via1 >>
rect 69 5694 121 5703
rect 69 5356 78 5694
rect 78 5356 112 5694
rect 112 5356 121 5694
rect 69 5347 121 5356
rect 15475 5694 15527 5703
rect 15475 5356 15484 5694
rect 15484 5356 15518 5694
rect 15518 5356 15527 5694
rect 15475 5347 15527 5356
rect 272 4708 324 4760
rect 572 4708 624 4760
rect 1172 4708 1224 4760
rect 1472 4708 1524 4760
rect 2072 4708 2124 4760
rect 2372 4708 2424 4760
rect 2972 4708 3024 4760
rect 3272 4708 3324 4760
rect 3872 4708 3924 4760
rect 4172 4708 4224 4760
rect 4772 4708 4824 4760
rect 5072 4708 5124 4760
rect 5672 4708 5724 4760
rect 5972 4708 6024 4760
rect 6572 4708 6624 4760
rect 6872 4708 6924 4760
rect 7472 4708 7524 4760
rect 7772 4708 7824 4760
rect 8372 4708 8424 4760
rect 8672 4708 8724 4760
rect 9272 4708 9324 4760
rect 9572 4708 9624 4760
rect 10172 4708 10224 4760
rect 10472 4708 10524 4760
rect 11072 4708 11124 4760
rect 11372 4708 11424 4760
rect 11972 4708 12024 4760
rect 12272 4708 12324 4760
rect 12872 4708 12924 4760
rect 13172 4708 13224 4760
rect 13772 4708 13824 4760
rect 14072 4708 14124 4760
rect 14672 4708 14724 4760
rect 14972 4708 15024 4760
rect 272 4615 324 4667
rect 14972 4615 15024 4667
rect 572 4490 624 4542
rect 1172 4490 1224 4542
rect 10600 4490 10652 4542
rect 1472 4413 1524 4465
rect 2072 4413 2124 4465
rect 11197 4413 11249 4465
rect 899 4332 959 4392
rect 2372 4336 2424 4388
rect 2972 4336 3024 4388
rect 9158 4336 9210 4388
rect 15007 4332 15067 4392
rect 3272 4259 3324 4311
rect 3872 4259 3924 4311
rect 9855 4259 9907 4311
rect 4172 4182 4224 4234
rect 4772 4182 4824 4234
rect 7916 4182 7968 4234
rect 5072 4105 5124 4157
rect 5672 4105 5724 4157
rect 8513 4105 8565 4157
rect 5972 4028 6024 4080
rect 6474 4028 6526 4080
rect 6572 4028 6624 4080
rect 6872 3951 6924 4003
rect 7171 3951 7223 4003
rect 7472 3951 7524 4003
rect 5132 3874 5184 3926
rect 7772 3874 7824 3926
rect 8372 3874 8424 3926
rect 5829 3797 5881 3849
rect 8672 3797 8724 3849
rect 9272 3797 9324 3849
rect 3790 3720 3842 3772
rect 9572 3720 9624 3772
rect 10172 3720 10224 3772
rect 4487 3643 4539 3695
rect 10472 3643 10524 3695
rect 11072 3643 11124 3695
rect 2448 3566 2500 3618
rect 11372 3566 11424 3618
rect 11972 3566 12024 3618
rect 3145 3489 3197 3541
rect 12272 3489 12324 3541
rect 12872 3489 12924 3541
rect 1106 3412 1158 3464
rect 13172 3412 13224 3464
rect 13772 3412 13824 3464
rect 1803 3335 1855 3387
rect 14072 3335 14124 3387
rect 14672 3335 14724 3387
<< metal2 >>
rect 63 5703 127 5709
rect 63 5347 69 5703
rect 121 5347 127 5703
rect 63 5341 127 5347
rect 15469 5703 15533 5709
rect 15469 5347 15475 5703
rect 15527 5347 15533 5703
rect 15469 5341 15533 5347
rect 65 4092 125 5341
rect 266 4708 272 4760
rect 324 4708 330 4760
rect 566 4708 572 4760
rect 624 4708 630 4760
rect 1166 4708 1172 4760
rect 1224 4708 1230 4760
rect 1466 4708 1472 4760
rect 1524 4708 1530 4760
rect 2066 4708 2072 4760
rect 2124 4708 2130 4760
rect 2366 4708 2372 4760
rect 2424 4708 2430 4760
rect 2966 4708 2972 4760
rect 3024 4708 3030 4760
rect 3266 4708 3272 4760
rect 3324 4708 3330 4760
rect 3866 4708 3872 4760
rect 3924 4708 3930 4760
rect 4166 4708 4172 4760
rect 4224 4708 4230 4760
rect 4766 4708 4772 4760
rect 4824 4708 4830 4760
rect 5066 4708 5072 4760
rect 5124 4708 5130 4760
rect 5666 4708 5672 4760
rect 5724 4708 5730 4760
rect 5966 4708 5972 4760
rect 6024 4708 6030 4760
rect 6566 4708 6572 4760
rect 6624 4708 6630 4760
rect 6866 4708 6872 4760
rect 6924 4708 6930 4760
rect 7466 4708 7472 4760
rect 7524 4708 7530 4760
rect 7766 4708 7772 4760
rect 7824 4708 7830 4760
rect 8366 4708 8372 4760
rect 8424 4708 8430 4760
rect 8666 4708 8672 4760
rect 8724 4708 8730 4760
rect 9266 4708 9272 4760
rect 9324 4708 9330 4760
rect 9566 4708 9572 4760
rect 9624 4708 9630 4760
rect 10166 4708 10172 4760
rect 10224 4708 10230 4760
rect 10466 4708 10472 4760
rect 10524 4708 10530 4760
rect 11066 4708 11072 4760
rect 11124 4708 11130 4760
rect 11366 4708 11372 4760
rect 11424 4708 11430 4760
rect 11966 4708 11972 4760
rect 12024 4708 12030 4760
rect 12266 4708 12272 4760
rect 12324 4708 12330 4760
rect 12866 4708 12872 4760
rect 12924 4708 12930 4760
rect 13166 4708 13172 4760
rect 13224 4708 13230 4760
rect 13766 4708 13772 4760
rect 13824 4708 13830 4760
rect 14066 4708 14072 4760
rect 14124 4708 14130 4760
rect 14666 4708 14672 4760
rect 14724 4708 14730 4760
rect 14966 4708 14972 4760
rect 15024 4708 15030 4760
rect 281 4667 315 4708
rect 266 4615 272 4667
rect 324 4615 330 4667
rect 581 4542 615 4708
rect 1181 4542 1215 4708
rect 566 4490 572 4542
rect 624 4490 630 4542
rect 1166 4490 1172 4542
rect 1224 4490 1230 4542
rect 1481 4465 1515 4708
rect 2081 4465 2115 4708
rect 1466 4413 1472 4465
rect 1524 4413 1530 4465
rect 2066 4413 2072 4465
rect 2124 4413 2130 4465
rect 893 4332 899 4392
rect 959 4332 965 4392
rect 2381 4388 2415 4708
rect 2981 4388 3015 4708
rect 2366 4336 2372 4388
rect 2424 4336 2430 4388
rect 2966 4336 2972 4388
rect 3024 4336 3030 4388
rect 65 4032 659 4092
rect 599 2972 659 4032
rect 592 2916 601 2972
rect 657 2916 666 2972
rect 599 2372 659 2916
rect 899 2672 959 4332
rect 3281 4311 3315 4708
rect 3881 4311 3915 4708
rect 3266 4259 3272 4311
rect 3324 4259 3330 4311
rect 3866 4259 3872 4311
rect 3924 4259 3930 4311
rect 4181 4234 4215 4708
rect 4781 4234 4815 4708
rect 4166 4182 4172 4234
rect 4224 4182 4230 4234
rect 4766 4182 4772 4234
rect 4824 4182 4830 4234
rect 5081 4157 5115 4708
rect 5681 4157 5715 4708
rect 5066 4105 5072 4157
rect 5124 4105 5130 4157
rect 5666 4105 5672 4157
rect 5724 4105 5730 4157
rect 5981 4080 6015 4708
rect 6581 4080 6615 4708
rect 5966 4028 5972 4080
rect 6024 4028 6030 4080
rect 6468 4028 6474 4080
rect 6526 4028 6532 4080
rect 6566 4028 6572 4080
rect 6624 4028 6630 4080
rect 5126 3874 5132 3926
rect 5184 3874 5190 3926
rect 3784 3720 3790 3772
rect 3842 3720 3848 3772
rect 2442 3566 2448 3618
rect 2500 3566 2506 3618
rect 1100 3412 1106 3464
rect 1158 3412 1164 3464
rect 1115 3189 1149 3412
rect 1797 3335 1803 3387
rect 1855 3335 1861 3387
rect 1812 3189 1846 3335
rect 2457 3189 2491 3566
rect 3139 3489 3145 3541
rect 3197 3489 3203 3541
rect 3154 3189 3188 3489
rect 3799 3189 3833 3720
rect 4481 3643 4487 3695
rect 4539 3643 4545 3695
rect 4496 3189 4530 3643
rect 5141 3189 5175 3874
rect 5823 3797 5829 3849
rect 5881 3797 5887 3849
rect 5838 3189 5872 3797
rect 6483 3189 6517 4028
rect 6881 4003 6915 4708
rect 7481 4003 7515 4708
rect 6866 3951 6872 4003
rect 6924 3951 6930 4003
rect 7165 3951 7171 4003
rect 7223 3951 7229 4003
rect 7466 3951 7472 4003
rect 7524 3951 7530 4003
rect 7180 3189 7214 3951
rect 7781 3926 7815 4708
rect 7910 4182 7916 4234
rect 7968 4182 7974 4234
rect 7766 3874 7772 3926
rect 7824 3874 7830 3926
rect 7925 3609 7959 4182
rect 8381 3926 8415 4708
rect 8507 4105 8513 4157
rect 8565 4105 8571 4157
rect 8366 3874 8372 3926
rect 8424 3874 8430 3926
rect 7825 3575 7959 3609
rect 7825 3189 7859 3575
rect 8522 3189 8556 4105
rect 8681 3849 8715 4708
rect 9152 4336 9158 4388
rect 9210 4336 9216 4388
rect 8666 3797 8672 3849
rect 8724 3797 8730 3849
rect 9167 3189 9201 4336
rect 9281 3849 9315 4708
rect 9266 3797 9272 3849
rect 9324 3797 9330 3849
rect 9581 3772 9615 4708
rect 9849 4259 9855 4311
rect 9907 4259 9913 4311
rect 9566 3720 9572 3772
rect 9624 3720 9630 3772
rect 9864 3189 9898 4259
rect 10181 3772 10215 4708
rect 10166 3720 10172 3772
rect 10224 3720 10230 3772
rect 10481 3695 10515 4708
rect 10594 4490 10600 4542
rect 10652 4490 10658 4542
rect 10466 3643 10472 3695
rect 10524 3643 10530 3695
rect 10609 3609 10643 4490
rect 11081 3695 11115 4708
rect 11191 4413 11197 4465
rect 11249 4413 11255 4465
rect 11066 3643 11072 3695
rect 11124 3643 11130 3695
rect 10509 3575 10643 3609
rect 10509 3189 10543 3575
rect 11206 3189 11240 4413
rect 11381 3618 11415 4708
rect 11981 3618 12015 4708
rect 11366 3566 11372 3618
rect 11424 3566 11430 3618
rect 11966 3566 11972 3618
rect 12024 3566 12030 3618
rect 12281 3541 12315 4708
rect 12881 3541 12915 4708
rect 12266 3489 12272 3541
rect 12324 3489 12330 3541
rect 12866 3489 12872 3541
rect 12924 3489 12930 3541
rect 13181 3464 13215 4708
rect 13781 3464 13815 4708
rect 13166 3412 13172 3464
rect 13224 3412 13230 3464
rect 13766 3412 13772 3464
rect 13824 3412 13830 3464
rect 14081 3387 14115 4708
rect 14681 3387 14715 4708
rect 14981 4667 15015 4708
rect 14966 4615 14972 4667
rect 15024 4615 15030 4667
rect 15001 4332 15007 4392
rect 15067 4332 15073 4392
rect 14066 3335 14072 3387
rect 14124 3335 14130 3387
rect 14666 3335 14672 3387
rect 14724 3335 14730 3387
rect 15007 2672 15067 4332
rect 15471 4092 15531 5341
rect 15307 4032 15531 4092
rect 15307 2972 15367 4032
rect 15300 2916 15309 2972
rect 15365 2916 15374 2972
rect 892 2616 901 2672
rect 957 2616 966 2672
rect 15000 2616 15009 2672
rect 15065 2616 15074 2672
rect 592 2316 601 2372
rect 657 2316 666 2372
rect 599 1772 659 2316
rect 899 2072 959 2616
rect 15007 2072 15067 2616
rect 15307 2372 15367 2916
rect 15300 2316 15309 2372
rect 15365 2316 15374 2372
rect 892 2016 901 2072
rect 957 2016 966 2072
rect 15000 2016 15009 2072
rect 15065 2016 15074 2072
rect 592 1716 601 1772
rect 657 1716 666 1772
rect 599 1172 659 1716
rect 899 1472 959 2016
rect 15007 1472 15067 2016
rect 15307 1772 15367 2316
rect 15300 1716 15309 1772
rect 15365 1716 15374 1772
rect 892 1416 901 1472
rect 957 1416 966 1472
rect 15000 1416 15009 1472
rect 15065 1416 15074 1472
rect 592 1116 601 1172
rect 657 1116 666 1172
rect 599 572 659 1116
rect 899 872 959 1416
rect 892 816 901 872
rect 957 816 966 872
rect 592 516 601 572
rect 657 516 666 572
rect 9864 0 9898 877
rect 11206 0 11240 877
rect 12548 0 12582 877
rect 13890 0 13924 877
rect 15007 872 15067 1416
rect 15307 1172 15367 1716
rect 15300 1116 15309 1172
rect 15365 1116 15374 1172
rect 15000 816 15009 872
rect 15065 816 15074 872
rect 15007 814 15067 816
rect 14236 572 14300 629
rect 15307 572 15367 1116
rect 14231 516 14240 572
rect 14296 516 14305 572
rect 15300 516 15309 572
rect 15365 516 15374 572
rect 14236 514 14300 516
rect 15307 514 15367 516
rect 14251 453 14285 514
<< via2 >>
rect 601 2916 657 2972
rect 15309 2916 15365 2972
rect 901 2616 957 2672
rect 15009 2616 15065 2672
rect 601 2316 657 2372
rect 15309 2316 15365 2372
rect 901 2016 957 2072
rect 15009 2016 15065 2072
rect 601 1716 657 1772
rect 15309 1716 15365 1772
rect 901 1416 957 1472
rect 15009 1416 15065 1472
rect 601 1116 657 1172
rect 901 816 957 872
rect 601 516 657 572
rect 15309 1116 15365 1172
rect 15009 816 15065 872
rect 14240 516 14296 572
rect 15309 516 15365 572
<< metal3 >>
rect 596 2974 662 2977
rect 15304 2974 15370 2977
rect 596 2972 15370 2974
rect 596 2916 601 2972
rect 657 2916 15309 2972
rect 15365 2916 15370 2972
rect 596 2914 15370 2916
rect 596 2911 662 2914
rect 15304 2911 15370 2914
rect 896 2674 962 2677
rect 15004 2674 15070 2677
rect 896 2672 15070 2674
rect 896 2616 901 2672
rect 957 2616 15009 2672
rect 15065 2616 15070 2672
rect 896 2614 15070 2616
rect 896 2611 962 2614
rect 15004 2611 15070 2614
rect 596 2374 662 2377
rect 15304 2374 15370 2377
rect 596 2372 15370 2374
rect 596 2316 601 2372
rect 657 2316 15309 2372
rect 15365 2316 15370 2372
rect 596 2314 15370 2316
rect 596 2311 662 2314
rect 15304 2311 15370 2314
rect 896 2074 962 2077
rect 15004 2074 15070 2077
rect 896 2072 15070 2074
rect 896 2016 901 2072
rect 957 2016 15009 2072
rect 15065 2016 15070 2072
rect 896 2014 15070 2016
rect 896 2011 962 2014
rect 15004 2011 15070 2014
rect 596 1774 662 1777
rect 15304 1774 15370 1777
rect 596 1772 15370 1774
rect 596 1716 601 1772
rect 657 1716 15309 1772
rect 15365 1716 15370 1772
rect 596 1714 15370 1716
rect 596 1711 662 1714
rect 15304 1711 15370 1714
rect 896 1474 962 1477
rect 15004 1474 15070 1477
rect 896 1472 15070 1474
rect 896 1416 901 1472
rect 957 1416 15009 1472
rect 15065 1416 15070 1472
rect 896 1414 15070 1416
rect 896 1411 962 1414
rect 15004 1411 15070 1414
rect 596 1174 662 1177
rect 15304 1174 15370 1177
rect 596 1172 15370 1174
rect 596 1116 601 1172
rect 657 1116 15309 1172
rect 15365 1116 15370 1172
rect 596 1114 15370 1116
rect 596 1111 662 1114
rect 15304 1111 15370 1114
rect 896 874 962 877
rect 15004 874 15070 877
rect 896 872 15070 874
rect 896 816 901 872
rect 957 816 15009 872
rect 15065 816 15070 872
rect 896 814 15070 816
rect 896 811 962 814
rect 15004 811 15070 814
rect 596 574 662 577
rect 14235 574 14301 577
rect 15304 574 15370 577
rect 596 572 15370 574
rect 596 516 601 572
rect 657 516 14240 572
rect 14296 516 15309 572
rect 15365 516 15370 572
rect 596 514 15370 516
rect 596 511 662 514
rect 14235 511 14301 514
rect 15304 511 15370 514
use decoder4  decoder4_0
timestamp 1748318706
transform 0 -1 14503 1 0 305
box -305 0 2996 13410
use shift_or2  shift_or2_0
timestamp 1748318706
transform 1 0 0 0 1 0
box 0 3329 15596 5868
<< labels >>
flabel metal1 15372 4785 15406 5629 1 FreeSans 128 0 0 0 C[16]
port 22 nsew signal output
flabel metal1 14472 4785 14506 5629 1 FreeSans 128 0 0 0 C[15]
port 21 nsew signal output
flabel metal1 13572 4785 13606 5629 1 FreeSans 128 0 0 0 C[14]
port 20 nsew signal output
flabel metal1 12672 4785 12706 5629 1 FreeSans 128 0 0 0 C[13]
port 19 nsew signal output
flabel metal1 11772 4785 11806 5629 1 FreeSans 128 0 0 0 C[12]
port 18 nsew signal output
flabel metal1 10872 4785 10906 5629 1 FreeSans 128 0 0 0 C[11]
port 17 nsew signal output
flabel metal1 9972 4785 10006 5629 1 FreeSans 128 0 0 0 C[10]
port 16 nsew signal output
flabel metal1 9072 4785 9106 5629 1 FreeSans 128 0 0 0 C[9]
port 15 nsew signal output
flabel metal1 8172 4785 8206 5629 1 FreeSans 128 0 0 0 C[8]
port 14 nsew signal output
flabel metal1 7272 4785 7306 5629 1 FreeSans 128 0 0 0 C[7]
port 13 nsew signal output
flabel metal1 6372 4785 6406 5629 1 FreeSans 128 0 0 0 C[6]
port 12 nsew signal output
flabel metal1 5472 4785 5506 5629 1 FreeSans 128 0 0 0 C[5]
port 11 nsew signal output
flabel metal1 4572 4785 4606 5629 1 FreeSans 128 0 0 0 C[4]
port 10 nsew signal output
flabel metal1 3672 4785 3706 5629 1 FreeSans 128 0 0 0 C[3]
port 9 nsew signal output
flabel metal1 2772 4785 2806 5629 1 FreeSans 128 0 0 0 C[2]
port 8 nsew signal output
flabel metal1 1872 4785 1906 5629 1 FreeSans 128 0 0 0 C[1]
port 7 nsew signal output
flabel metal1 972 4785 1006 5629 1 FreeSans 128 0 0 0 C[0]
port 6 nsew signal output
flabel metal2 9864 0 9898 877 0 FreeSans 128 270 0 0 IN[5]
port 3 nsew signal input
flabel metal2 11206 0 11240 877 0 FreeSans 128 270 0 0 IN[4]
port 2 nsew signal input
flabel metal2 12548 0 12582 877 0 FreeSans 128 270 0 0 IN[7]
port 5 nsew signal input
flabel metal2 13890 0 13924 877 0 FreeSans 128 270 0 0 IN[6]
port 4 nsew signal input
flabel metal3 1199 814 14467 874 0 FreeSans 128 270 0 0 VSS
port 0 nsew ground bidirectional
flabel metal3 1199 514 14467 574 0 FreeSans 128 270 0 0 VDD
port 1 nsew power bidirectional
<< end >>
