magic
tech sky130A
magscale 1 2
timestamp 1748065934
<< nwell >>
rect -60 606 15536 1292
<< pwell >>
rect -60 556 126 557
rect -60 0 15536 556
<< mvnmos >>
rect 188 213 288 343
rect 488 213 588 343
rect 788 213 888 343
rect 1088 213 1188 343
rect 1388 213 1488 343
rect 1688 213 1788 343
rect 1988 213 2088 343
rect 2288 213 2388 343
rect 2588 213 2688 343
rect 2888 213 2988 343
rect 3188 213 3288 343
rect 3488 213 3588 343
rect 3788 213 3888 343
rect 4088 213 4188 343
rect 4388 213 4488 343
rect 4688 213 4788 343
rect 4988 213 5088 343
rect 5288 213 5388 343
rect 5588 213 5688 343
rect 5888 213 5988 343
rect 6188 213 6288 343
rect 6488 213 6588 343
rect 6788 213 6888 343
rect 7088 213 7188 343
rect 7388 213 7488 343
rect 7688 213 7788 343
rect 7988 213 8088 343
rect 8288 213 8388 343
rect 8588 213 8688 343
rect 8888 213 8988 343
rect 9188 213 9288 343
rect 9488 213 9588 343
rect 9788 213 9888 343
rect 10088 213 10188 343
rect 10388 213 10488 343
rect 10688 213 10788 343
rect 10988 213 11088 343
rect 11288 213 11388 343
rect 11588 213 11688 343
rect 11888 213 11988 343
rect 12188 213 12288 343
rect 12488 213 12588 343
rect 12788 213 12888 343
rect 13088 213 13188 343
rect 13388 213 13488 343
rect 13688 213 13788 343
rect 13988 213 14088 343
rect 14288 213 14388 343
rect 14588 213 14688 343
rect 14888 213 14988 343
rect 15188 213 15288 343
<< mvpmos >>
rect 188 849 288 1049
rect 488 849 588 1049
rect 788 849 888 1049
rect 1088 849 1188 1049
rect 1388 849 1488 1049
rect 1688 849 1788 1049
rect 1988 849 2088 1049
rect 2288 849 2388 1049
rect 2588 849 2688 1049
rect 2888 849 2988 1049
rect 3188 849 3288 1049
rect 3488 849 3588 1049
rect 3788 849 3888 1049
rect 4088 849 4188 1049
rect 4388 849 4488 1049
rect 4688 849 4788 1049
rect 4988 849 5088 1049
rect 5288 849 5388 1049
rect 5588 849 5688 1049
rect 5888 849 5988 1049
rect 6188 849 6288 1049
rect 6488 849 6588 1049
rect 6788 849 6888 1049
rect 7088 849 7188 1049
rect 7388 849 7488 1049
rect 7688 849 7788 1049
rect 7988 849 8088 1049
rect 8288 849 8388 1049
rect 8588 849 8688 1049
rect 8888 849 8988 1049
rect 9188 849 9288 1049
rect 9488 849 9588 1049
rect 9788 849 9888 1049
rect 10088 849 10188 1049
rect 10388 849 10488 1049
rect 10688 849 10788 1049
rect 10988 849 11088 1049
rect 11288 849 11388 1049
rect 11588 849 11688 1049
rect 11888 849 11988 1049
rect 12188 849 12288 1049
rect 12488 849 12588 1049
rect 12788 849 12888 1049
rect 13088 849 13188 1049
rect 13388 849 13488 1049
rect 13688 849 13788 1049
rect 13988 849 14088 1049
rect 14288 849 14388 1049
rect 14588 849 14688 1049
rect 14888 849 14988 1049
rect 15188 849 15288 1049
<< mvndiff >>
rect 118 331 188 343
rect 118 225 130 331
rect 164 225 188 331
rect 118 213 188 225
rect 288 331 358 343
rect 288 225 312 331
rect 346 225 358 331
rect 288 213 358 225
rect 418 331 488 343
rect 418 225 430 331
rect 464 225 488 331
rect 418 213 488 225
rect 588 331 658 343
rect 588 225 612 331
rect 646 225 658 331
rect 588 213 658 225
rect 718 331 788 343
rect 718 225 730 331
rect 764 225 788 331
rect 718 213 788 225
rect 888 331 958 343
rect 888 225 912 331
rect 946 225 958 331
rect 888 213 958 225
rect 1018 331 1088 343
rect 1018 225 1030 331
rect 1064 225 1088 331
rect 1018 213 1088 225
rect 1188 331 1258 343
rect 1188 225 1212 331
rect 1246 225 1258 331
rect 1188 213 1258 225
rect 1318 331 1388 343
rect 1318 225 1330 331
rect 1364 225 1388 331
rect 1318 213 1388 225
rect 1488 331 1558 343
rect 1488 225 1512 331
rect 1546 225 1558 331
rect 1488 213 1558 225
rect 1618 331 1688 343
rect 1618 225 1630 331
rect 1664 225 1688 331
rect 1618 213 1688 225
rect 1788 331 1858 343
rect 1788 225 1812 331
rect 1846 225 1858 331
rect 1788 213 1858 225
rect 1918 331 1988 343
rect 1918 225 1930 331
rect 1964 225 1988 331
rect 1918 213 1988 225
rect 2088 331 2158 343
rect 2088 225 2112 331
rect 2146 225 2158 331
rect 2088 213 2158 225
rect 2218 331 2288 343
rect 2218 225 2230 331
rect 2264 225 2288 331
rect 2218 213 2288 225
rect 2388 331 2458 343
rect 2388 225 2412 331
rect 2446 225 2458 331
rect 2388 213 2458 225
rect 2518 331 2588 343
rect 2518 225 2530 331
rect 2564 225 2588 331
rect 2518 213 2588 225
rect 2688 331 2758 343
rect 2688 225 2712 331
rect 2746 225 2758 331
rect 2688 213 2758 225
rect 2818 331 2888 343
rect 2818 225 2830 331
rect 2864 225 2888 331
rect 2818 213 2888 225
rect 2988 331 3058 343
rect 2988 225 3012 331
rect 3046 225 3058 331
rect 2988 213 3058 225
rect 3118 331 3188 343
rect 3118 225 3130 331
rect 3164 225 3188 331
rect 3118 213 3188 225
rect 3288 331 3358 343
rect 3288 225 3312 331
rect 3346 225 3358 331
rect 3288 213 3358 225
rect 3418 331 3488 343
rect 3418 225 3430 331
rect 3464 225 3488 331
rect 3418 213 3488 225
rect 3588 331 3658 343
rect 3588 225 3612 331
rect 3646 225 3658 331
rect 3588 213 3658 225
rect 3718 331 3788 343
rect 3718 225 3730 331
rect 3764 225 3788 331
rect 3718 213 3788 225
rect 3888 331 3958 343
rect 3888 225 3912 331
rect 3946 225 3958 331
rect 3888 213 3958 225
rect 4018 331 4088 343
rect 4018 225 4030 331
rect 4064 225 4088 331
rect 4018 213 4088 225
rect 4188 331 4258 343
rect 4188 225 4212 331
rect 4246 225 4258 331
rect 4188 213 4258 225
rect 4318 331 4388 343
rect 4318 225 4330 331
rect 4364 225 4388 331
rect 4318 213 4388 225
rect 4488 331 4558 343
rect 4488 225 4512 331
rect 4546 225 4558 331
rect 4488 213 4558 225
rect 4618 331 4688 343
rect 4618 225 4630 331
rect 4664 225 4688 331
rect 4618 213 4688 225
rect 4788 331 4858 343
rect 4788 225 4812 331
rect 4846 225 4858 331
rect 4788 213 4858 225
rect 4918 331 4988 343
rect 4918 225 4930 331
rect 4964 225 4988 331
rect 4918 213 4988 225
rect 5088 331 5158 343
rect 5088 225 5112 331
rect 5146 225 5158 331
rect 5088 213 5158 225
rect 5218 331 5288 343
rect 5218 225 5230 331
rect 5264 225 5288 331
rect 5218 213 5288 225
rect 5388 331 5458 343
rect 5388 225 5412 331
rect 5446 225 5458 331
rect 5388 213 5458 225
rect 5518 331 5588 343
rect 5518 225 5530 331
rect 5564 225 5588 331
rect 5518 213 5588 225
rect 5688 331 5758 343
rect 5688 225 5712 331
rect 5746 225 5758 331
rect 5688 213 5758 225
rect 5818 331 5888 343
rect 5818 225 5830 331
rect 5864 225 5888 331
rect 5818 213 5888 225
rect 5988 331 6058 343
rect 5988 225 6012 331
rect 6046 225 6058 331
rect 5988 213 6058 225
rect 6118 331 6188 343
rect 6118 225 6130 331
rect 6164 225 6188 331
rect 6118 213 6188 225
rect 6288 331 6358 343
rect 6288 225 6312 331
rect 6346 225 6358 331
rect 6288 213 6358 225
rect 6418 331 6488 343
rect 6418 225 6430 331
rect 6464 225 6488 331
rect 6418 213 6488 225
rect 6588 331 6658 343
rect 6588 225 6612 331
rect 6646 225 6658 331
rect 6588 213 6658 225
rect 6718 331 6788 343
rect 6718 225 6730 331
rect 6764 225 6788 331
rect 6718 213 6788 225
rect 6888 331 6958 343
rect 6888 225 6912 331
rect 6946 225 6958 331
rect 6888 213 6958 225
rect 7018 331 7088 343
rect 7018 225 7030 331
rect 7064 225 7088 331
rect 7018 213 7088 225
rect 7188 331 7258 343
rect 7188 225 7212 331
rect 7246 225 7258 331
rect 7188 213 7258 225
rect 7318 331 7388 343
rect 7318 225 7330 331
rect 7364 225 7388 331
rect 7318 213 7388 225
rect 7488 331 7558 343
rect 7488 225 7512 331
rect 7546 225 7558 331
rect 7488 213 7558 225
rect 7618 331 7688 343
rect 7618 225 7630 331
rect 7664 225 7688 331
rect 7618 213 7688 225
rect 7788 331 7858 343
rect 7788 225 7812 331
rect 7846 225 7858 331
rect 7788 213 7858 225
rect 7918 331 7988 343
rect 7918 225 7930 331
rect 7964 225 7988 331
rect 7918 213 7988 225
rect 8088 331 8158 343
rect 8088 225 8112 331
rect 8146 225 8158 331
rect 8088 213 8158 225
rect 8218 331 8288 343
rect 8218 225 8230 331
rect 8264 225 8288 331
rect 8218 213 8288 225
rect 8388 331 8458 343
rect 8388 225 8412 331
rect 8446 225 8458 331
rect 8388 213 8458 225
rect 8518 331 8588 343
rect 8518 225 8530 331
rect 8564 225 8588 331
rect 8518 213 8588 225
rect 8688 331 8758 343
rect 8688 225 8712 331
rect 8746 225 8758 331
rect 8688 213 8758 225
rect 8818 331 8888 343
rect 8818 225 8830 331
rect 8864 225 8888 331
rect 8818 213 8888 225
rect 8988 331 9058 343
rect 8988 225 9012 331
rect 9046 225 9058 331
rect 8988 213 9058 225
rect 9118 331 9188 343
rect 9118 225 9130 331
rect 9164 225 9188 331
rect 9118 213 9188 225
rect 9288 331 9358 343
rect 9288 225 9312 331
rect 9346 225 9358 331
rect 9288 213 9358 225
rect 9418 331 9488 343
rect 9418 225 9430 331
rect 9464 225 9488 331
rect 9418 213 9488 225
rect 9588 331 9658 343
rect 9588 225 9612 331
rect 9646 225 9658 331
rect 9588 213 9658 225
rect 9718 331 9788 343
rect 9718 225 9730 331
rect 9764 225 9788 331
rect 9718 213 9788 225
rect 9888 331 9958 343
rect 9888 225 9912 331
rect 9946 225 9958 331
rect 9888 213 9958 225
rect 10018 331 10088 343
rect 10018 225 10030 331
rect 10064 225 10088 331
rect 10018 213 10088 225
rect 10188 331 10258 343
rect 10188 225 10212 331
rect 10246 225 10258 331
rect 10188 213 10258 225
rect 10318 331 10388 343
rect 10318 225 10330 331
rect 10364 225 10388 331
rect 10318 213 10388 225
rect 10488 331 10558 343
rect 10488 225 10512 331
rect 10546 225 10558 331
rect 10488 213 10558 225
rect 10618 331 10688 343
rect 10618 225 10630 331
rect 10664 225 10688 331
rect 10618 213 10688 225
rect 10788 331 10858 343
rect 10788 225 10812 331
rect 10846 225 10858 331
rect 10788 213 10858 225
rect 10918 331 10988 343
rect 10918 225 10930 331
rect 10964 225 10988 331
rect 10918 213 10988 225
rect 11088 331 11158 343
rect 11088 225 11112 331
rect 11146 225 11158 331
rect 11088 213 11158 225
rect 11218 331 11288 343
rect 11218 225 11230 331
rect 11264 225 11288 331
rect 11218 213 11288 225
rect 11388 331 11458 343
rect 11388 225 11412 331
rect 11446 225 11458 331
rect 11388 213 11458 225
rect 11518 331 11588 343
rect 11518 225 11530 331
rect 11564 225 11588 331
rect 11518 213 11588 225
rect 11688 331 11758 343
rect 11688 225 11712 331
rect 11746 225 11758 331
rect 11688 213 11758 225
rect 11818 331 11888 343
rect 11818 225 11830 331
rect 11864 225 11888 331
rect 11818 213 11888 225
rect 11988 331 12058 343
rect 11988 225 12012 331
rect 12046 225 12058 331
rect 11988 213 12058 225
rect 12118 331 12188 343
rect 12118 225 12130 331
rect 12164 225 12188 331
rect 12118 213 12188 225
rect 12288 331 12358 343
rect 12288 225 12312 331
rect 12346 225 12358 331
rect 12288 213 12358 225
rect 12418 331 12488 343
rect 12418 225 12430 331
rect 12464 225 12488 331
rect 12418 213 12488 225
rect 12588 331 12658 343
rect 12588 225 12612 331
rect 12646 225 12658 331
rect 12588 213 12658 225
rect 12718 331 12788 343
rect 12718 225 12730 331
rect 12764 225 12788 331
rect 12718 213 12788 225
rect 12888 331 12958 343
rect 12888 225 12912 331
rect 12946 225 12958 331
rect 12888 213 12958 225
rect 13018 331 13088 343
rect 13018 225 13030 331
rect 13064 225 13088 331
rect 13018 213 13088 225
rect 13188 331 13258 343
rect 13188 225 13212 331
rect 13246 225 13258 331
rect 13188 213 13258 225
rect 13318 331 13388 343
rect 13318 225 13330 331
rect 13364 225 13388 331
rect 13318 213 13388 225
rect 13488 331 13558 343
rect 13488 225 13512 331
rect 13546 225 13558 331
rect 13488 213 13558 225
rect 13618 331 13688 343
rect 13618 225 13630 331
rect 13664 225 13688 331
rect 13618 213 13688 225
rect 13788 331 13858 343
rect 13788 225 13812 331
rect 13846 225 13858 331
rect 13788 213 13858 225
rect 13918 331 13988 343
rect 13918 225 13930 331
rect 13964 225 13988 331
rect 13918 213 13988 225
rect 14088 331 14158 343
rect 14088 225 14112 331
rect 14146 225 14158 331
rect 14088 213 14158 225
rect 14218 331 14288 343
rect 14218 225 14230 331
rect 14264 225 14288 331
rect 14218 213 14288 225
rect 14388 331 14458 343
rect 14388 225 14412 331
rect 14446 225 14458 331
rect 14388 213 14458 225
rect 14518 331 14588 343
rect 14518 225 14530 331
rect 14564 225 14588 331
rect 14518 213 14588 225
rect 14688 331 14758 343
rect 14688 225 14712 331
rect 14746 225 14758 331
rect 14688 213 14758 225
rect 14818 331 14888 343
rect 14818 225 14830 331
rect 14864 225 14888 331
rect 14818 213 14888 225
rect 14988 331 15058 343
rect 14988 225 15012 331
rect 15046 225 15058 331
rect 14988 213 15058 225
rect 15118 331 15188 343
rect 15118 225 15130 331
rect 15164 225 15188 331
rect 15118 213 15188 225
rect 15288 331 15358 343
rect 15288 225 15312 331
rect 15346 225 15358 331
rect 15288 213 15358 225
<< mvpdiff >>
rect 118 1037 188 1049
rect 118 861 130 1037
rect 164 861 188 1037
rect 118 849 188 861
rect 288 1037 358 1049
rect 288 861 312 1037
rect 346 861 358 1037
rect 288 849 358 861
rect 418 1037 488 1049
rect 418 861 430 1037
rect 464 861 488 1037
rect 418 849 488 861
rect 588 1037 658 1049
rect 588 861 612 1037
rect 646 861 658 1037
rect 588 849 658 861
rect 718 1037 788 1049
rect 718 861 730 1037
rect 764 861 788 1037
rect 718 849 788 861
rect 888 1037 958 1049
rect 888 861 912 1037
rect 946 861 958 1037
rect 888 849 958 861
rect 1018 1037 1088 1049
rect 1018 861 1030 1037
rect 1064 861 1088 1037
rect 1018 849 1088 861
rect 1188 1037 1258 1049
rect 1188 861 1212 1037
rect 1246 861 1258 1037
rect 1188 849 1258 861
rect 1318 1037 1388 1049
rect 1318 861 1330 1037
rect 1364 861 1388 1037
rect 1318 849 1388 861
rect 1488 1037 1558 1049
rect 1488 861 1512 1037
rect 1546 861 1558 1037
rect 1488 849 1558 861
rect 1618 1037 1688 1049
rect 1618 861 1630 1037
rect 1664 861 1688 1037
rect 1618 849 1688 861
rect 1788 1037 1858 1049
rect 1788 861 1812 1037
rect 1846 861 1858 1037
rect 1788 849 1858 861
rect 1918 1037 1988 1049
rect 1918 861 1930 1037
rect 1964 861 1988 1037
rect 1918 849 1988 861
rect 2088 1037 2158 1049
rect 2088 861 2112 1037
rect 2146 861 2158 1037
rect 2088 849 2158 861
rect 2218 1037 2288 1049
rect 2218 861 2230 1037
rect 2264 861 2288 1037
rect 2218 849 2288 861
rect 2388 1037 2458 1049
rect 2388 861 2412 1037
rect 2446 861 2458 1037
rect 2388 849 2458 861
rect 2518 1037 2588 1049
rect 2518 861 2530 1037
rect 2564 861 2588 1037
rect 2518 849 2588 861
rect 2688 1037 2758 1049
rect 2688 861 2712 1037
rect 2746 861 2758 1037
rect 2688 849 2758 861
rect 2818 1037 2888 1049
rect 2818 861 2830 1037
rect 2864 861 2888 1037
rect 2818 849 2888 861
rect 2988 1037 3058 1049
rect 2988 861 3012 1037
rect 3046 861 3058 1037
rect 2988 849 3058 861
rect 3118 1037 3188 1049
rect 3118 861 3130 1037
rect 3164 861 3188 1037
rect 3118 849 3188 861
rect 3288 1037 3358 1049
rect 3288 861 3312 1037
rect 3346 861 3358 1037
rect 3288 849 3358 861
rect 3418 1037 3488 1049
rect 3418 861 3430 1037
rect 3464 861 3488 1037
rect 3418 849 3488 861
rect 3588 1037 3658 1049
rect 3588 861 3612 1037
rect 3646 861 3658 1037
rect 3588 849 3658 861
rect 3718 1037 3788 1049
rect 3718 861 3730 1037
rect 3764 861 3788 1037
rect 3718 849 3788 861
rect 3888 1037 3958 1049
rect 3888 861 3912 1037
rect 3946 861 3958 1037
rect 3888 849 3958 861
rect 4018 1037 4088 1049
rect 4018 861 4030 1037
rect 4064 861 4088 1037
rect 4018 849 4088 861
rect 4188 1037 4258 1049
rect 4188 861 4212 1037
rect 4246 861 4258 1037
rect 4188 849 4258 861
rect 4318 1037 4388 1049
rect 4318 861 4330 1037
rect 4364 861 4388 1037
rect 4318 849 4388 861
rect 4488 1037 4558 1049
rect 4488 861 4512 1037
rect 4546 861 4558 1037
rect 4488 849 4558 861
rect 4618 1037 4688 1049
rect 4618 861 4630 1037
rect 4664 861 4688 1037
rect 4618 849 4688 861
rect 4788 1037 4858 1049
rect 4788 861 4812 1037
rect 4846 861 4858 1037
rect 4788 849 4858 861
rect 4918 1037 4988 1049
rect 4918 861 4930 1037
rect 4964 861 4988 1037
rect 4918 849 4988 861
rect 5088 1037 5158 1049
rect 5088 861 5112 1037
rect 5146 861 5158 1037
rect 5088 849 5158 861
rect 5218 1037 5288 1049
rect 5218 861 5230 1037
rect 5264 861 5288 1037
rect 5218 849 5288 861
rect 5388 1037 5458 1049
rect 5388 861 5412 1037
rect 5446 861 5458 1037
rect 5388 849 5458 861
rect 5518 1037 5588 1049
rect 5518 861 5530 1037
rect 5564 861 5588 1037
rect 5518 849 5588 861
rect 5688 1037 5758 1049
rect 5688 861 5712 1037
rect 5746 861 5758 1037
rect 5688 849 5758 861
rect 5818 1037 5888 1049
rect 5818 861 5830 1037
rect 5864 861 5888 1037
rect 5818 849 5888 861
rect 5988 1037 6058 1049
rect 5988 861 6012 1037
rect 6046 861 6058 1037
rect 5988 849 6058 861
rect 6118 1037 6188 1049
rect 6118 861 6130 1037
rect 6164 861 6188 1037
rect 6118 849 6188 861
rect 6288 1037 6358 1049
rect 6288 861 6312 1037
rect 6346 861 6358 1037
rect 6288 849 6358 861
rect 6418 1037 6488 1049
rect 6418 861 6430 1037
rect 6464 861 6488 1037
rect 6418 849 6488 861
rect 6588 1037 6658 1049
rect 6588 861 6612 1037
rect 6646 861 6658 1037
rect 6588 849 6658 861
rect 6718 1037 6788 1049
rect 6718 861 6730 1037
rect 6764 861 6788 1037
rect 6718 849 6788 861
rect 6888 1037 6958 1049
rect 6888 861 6912 1037
rect 6946 861 6958 1037
rect 6888 849 6958 861
rect 7018 1037 7088 1049
rect 7018 861 7030 1037
rect 7064 861 7088 1037
rect 7018 849 7088 861
rect 7188 1037 7258 1049
rect 7188 861 7212 1037
rect 7246 861 7258 1037
rect 7188 849 7258 861
rect 7318 1037 7388 1049
rect 7318 861 7330 1037
rect 7364 861 7388 1037
rect 7318 849 7388 861
rect 7488 1037 7558 1049
rect 7488 861 7512 1037
rect 7546 861 7558 1037
rect 7488 849 7558 861
rect 7618 1037 7688 1049
rect 7618 861 7630 1037
rect 7664 861 7688 1037
rect 7618 849 7688 861
rect 7788 1037 7858 1049
rect 7788 861 7812 1037
rect 7846 861 7858 1037
rect 7788 849 7858 861
rect 7918 1037 7988 1049
rect 7918 861 7930 1037
rect 7964 861 7988 1037
rect 7918 849 7988 861
rect 8088 1037 8158 1049
rect 8088 861 8112 1037
rect 8146 861 8158 1037
rect 8088 849 8158 861
rect 8218 1037 8288 1049
rect 8218 861 8230 1037
rect 8264 861 8288 1037
rect 8218 849 8288 861
rect 8388 1037 8458 1049
rect 8388 861 8412 1037
rect 8446 861 8458 1037
rect 8388 849 8458 861
rect 8518 1037 8588 1049
rect 8518 861 8530 1037
rect 8564 861 8588 1037
rect 8518 849 8588 861
rect 8688 1037 8758 1049
rect 8688 861 8712 1037
rect 8746 861 8758 1037
rect 8688 849 8758 861
rect 8818 1037 8888 1049
rect 8818 861 8830 1037
rect 8864 861 8888 1037
rect 8818 849 8888 861
rect 8988 1037 9058 1049
rect 8988 861 9012 1037
rect 9046 861 9058 1037
rect 8988 849 9058 861
rect 9118 1037 9188 1049
rect 9118 861 9130 1037
rect 9164 861 9188 1037
rect 9118 849 9188 861
rect 9288 1037 9358 1049
rect 9288 861 9312 1037
rect 9346 861 9358 1037
rect 9288 849 9358 861
rect 9418 1037 9488 1049
rect 9418 861 9430 1037
rect 9464 861 9488 1037
rect 9418 849 9488 861
rect 9588 1037 9658 1049
rect 9588 861 9612 1037
rect 9646 861 9658 1037
rect 9588 849 9658 861
rect 9718 1037 9788 1049
rect 9718 861 9730 1037
rect 9764 861 9788 1037
rect 9718 849 9788 861
rect 9888 1037 9958 1049
rect 9888 861 9912 1037
rect 9946 861 9958 1037
rect 9888 849 9958 861
rect 10018 1037 10088 1049
rect 10018 861 10030 1037
rect 10064 861 10088 1037
rect 10018 849 10088 861
rect 10188 1037 10258 1049
rect 10188 861 10212 1037
rect 10246 861 10258 1037
rect 10188 849 10258 861
rect 10318 1037 10388 1049
rect 10318 861 10330 1037
rect 10364 861 10388 1037
rect 10318 849 10388 861
rect 10488 1037 10558 1049
rect 10488 861 10512 1037
rect 10546 861 10558 1037
rect 10488 849 10558 861
rect 10618 1037 10688 1049
rect 10618 861 10630 1037
rect 10664 861 10688 1037
rect 10618 849 10688 861
rect 10788 1037 10858 1049
rect 10788 861 10812 1037
rect 10846 861 10858 1037
rect 10788 849 10858 861
rect 10918 1037 10988 1049
rect 10918 861 10930 1037
rect 10964 861 10988 1037
rect 10918 849 10988 861
rect 11088 1037 11158 1049
rect 11088 861 11112 1037
rect 11146 861 11158 1037
rect 11088 849 11158 861
rect 11218 1037 11288 1049
rect 11218 861 11230 1037
rect 11264 861 11288 1037
rect 11218 849 11288 861
rect 11388 1037 11458 1049
rect 11388 861 11412 1037
rect 11446 861 11458 1037
rect 11388 849 11458 861
rect 11518 1037 11588 1049
rect 11518 861 11530 1037
rect 11564 861 11588 1037
rect 11518 849 11588 861
rect 11688 1037 11758 1049
rect 11688 861 11712 1037
rect 11746 861 11758 1037
rect 11688 849 11758 861
rect 11818 1037 11888 1049
rect 11818 861 11830 1037
rect 11864 861 11888 1037
rect 11818 849 11888 861
rect 11988 1037 12058 1049
rect 11988 861 12012 1037
rect 12046 861 12058 1037
rect 11988 849 12058 861
rect 12118 1037 12188 1049
rect 12118 861 12130 1037
rect 12164 861 12188 1037
rect 12118 849 12188 861
rect 12288 1037 12358 1049
rect 12288 861 12312 1037
rect 12346 861 12358 1037
rect 12288 849 12358 861
rect 12418 1037 12488 1049
rect 12418 861 12430 1037
rect 12464 861 12488 1037
rect 12418 849 12488 861
rect 12588 1037 12658 1049
rect 12588 861 12612 1037
rect 12646 861 12658 1037
rect 12588 849 12658 861
rect 12718 1037 12788 1049
rect 12718 861 12730 1037
rect 12764 861 12788 1037
rect 12718 849 12788 861
rect 12888 1037 12958 1049
rect 12888 861 12912 1037
rect 12946 861 12958 1037
rect 12888 849 12958 861
rect 13018 1037 13088 1049
rect 13018 861 13030 1037
rect 13064 861 13088 1037
rect 13018 849 13088 861
rect 13188 1037 13258 1049
rect 13188 861 13212 1037
rect 13246 861 13258 1037
rect 13188 849 13258 861
rect 13318 1037 13388 1049
rect 13318 861 13330 1037
rect 13364 861 13388 1037
rect 13318 849 13388 861
rect 13488 1037 13558 1049
rect 13488 861 13512 1037
rect 13546 861 13558 1037
rect 13488 849 13558 861
rect 13618 1037 13688 1049
rect 13618 861 13630 1037
rect 13664 861 13688 1037
rect 13618 849 13688 861
rect 13788 1037 13858 1049
rect 13788 861 13812 1037
rect 13846 861 13858 1037
rect 13788 849 13858 861
rect 13918 1037 13988 1049
rect 13918 861 13930 1037
rect 13964 861 13988 1037
rect 13918 849 13988 861
rect 14088 1037 14158 1049
rect 14088 861 14112 1037
rect 14146 861 14158 1037
rect 14088 849 14158 861
rect 14218 1037 14288 1049
rect 14218 861 14230 1037
rect 14264 861 14288 1037
rect 14218 849 14288 861
rect 14388 1037 14458 1049
rect 14388 861 14412 1037
rect 14446 861 14458 1037
rect 14388 849 14458 861
rect 14518 1037 14588 1049
rect 14518 861 14530 1037
rect 14564 861 14588 1037
rect 14518 849 14588 861
rect 14688 1037 14758 1049
rect 14688 861 14712 1037
rect 14746 861 14758 1037
rect 14688 849 14758 861
rect 14818 1037 14888 1049
rect 14818 861 14830 1037
rect 14864 861 14888 1037
rect 14818 849 14888 861
rect 14988 1037 15058 1049
rect 14988 861 15012 1037
rect 15046 861 15058 1037
rect 14988 849 15058 861
rect 15118 1037 15188 1049
rect 15118 861 15130 1037
rect 15164 861 15188 1037
rect 15118 849 15188 861
rect 15288 1037 15358 1049
rect 15288 861 15312 1037
rect 15346 861 15358 1037
rect 15288 849 15358 861
<< mvndiffc >>
rect 130 225 164 331
rect 312 225 346 331
rect 430 225 464 331
rect 612 225 646 331
rect 730 225 764 331
rect 912 225 946 331
rect 1030 225 1064 331
rect 1212 225 1246 331
rect 1330 225 1364 331
rect 1512 225 1546 331
rect 1630 225 1664 331
rect 1812 225 1846 331
rect 1930 225 1964 331
rect 2112 225 2146 331
rect 2230 225 2264 331
rect 2412 225 2446 331
rect 2530 225 2564 331
rect 2712 225 2746 331
rect 2830 225 2864 331
rect 3012 225 3046 331
rect 3130 225 3164 331
rect 3312 225 3346 331
rect 3430 225 3464 331
rect 3612 225 3646 331
rect 3730 225 3764 331
rect 3912 225 3946 331
rect 4030 225 4064 331
rect 4212 225 4246 331
rect 4330 225 4364 331
rect 4512 225 4546 331
rect 4630 225 4664 331
rect 4812 225 4846 331
rect 4930 225 4964 331
rect 5112 225 5146 331
rect 5230 225 5264 331
rect 5412 225 5446 331
rect 5530 225 5564 331
rect 5712 225 5746 331
rect 5830 225 5864 331
rect 6012 225 6046 331
rect 6130 225 6164 331
rect 6312 225 6346 331
rect 6430 225 6464 331
rect 6612 225 6646 331
rect 6730 225 6764 331
rect 6912 225 6946 331
rect 7030 225 7064 331
rect 7212 225 7246 331
rect 7330 225 7364 331
rect 7512 225 7546 331
rect 7630 225 7664 331
rect 7812 225 7846 331
rect 7930 225 7964 331
rect 8112 225 8146 331
rect 8230 225 8264 331
rect 8412 225 8446 331
rect 8530 225 8564 331
rect 8712 225 8746 331
rect 8830 225 8864 331
rect 9012 225 9046 331
rect 9130 225 9164 331
rect 9312 225 9346 331
rect 9430 225 9464 331
rect 9612 225 9646 331
rect 9730 225 9764 331
rect 9912 225 9946 331
rect 10030 225 10064 331
rect 10212 225 10246 331
rect 10330 225 10364 331
rect 10512 225 10546 331
rect 10630 225 10664 331
rect 10812 225 10846 331
rect 10930 225 10964 331
rect 11112 225 11146 331
rect 11230 225 11264 331
rect 11412 225 11446 331
rect 11530 225 11564 331
rect 11712 225 11746 331
rect 11830 225 11864 331
rect 12012 225 12046 331
rect 12130 225 12164 331
rect 12312 225 12346 331
rect 12430 225 12464 331
rect 12612 225 12646 331
rect 12730 225 12764 331
rect 12912 225 12946 331
rect 13030 225 13064 331
rect 13212 225 13246 331
rect 13330 225 13364 331
rect 13512 225 13546 331
rect 13630 225 13664 331
rect 13812 225 13846 331
rect 13930 225 13964 331
rect 14112 225 14146 331
rect 14230 225 14264 331
rect 14412 225 14446 331
rect 14530 225 14564 331
rect 14712 225 14746 331
rect 14830 225 14864 331
rect 15012 225 15046 331
rect 15130 225 15164 331
rect 15312 225 15346 331
<< mvpdiffc >>
rect 130 861 164 1037
rect 312 861 346 1037
rect 430 861 464 1037
rect 612 861 646 1037
rect 730 861 764 1037
rect 912 861 946 1037
rect 1030 861 1064 1037
rect 1212 861 1246 1037
rect 1330 861 1364 1037
rect 1512 861 1546 1037
rect 1630 861 1664 1037
rect 1812 861 1846 1037
rect 1930 861 1964 1037
rect 2112 861 2146 1037
rect 2230 861 2264 1037
rect 2412 861 2446 1037
rect 2530 861 2564 1037
rect 2712 861 2746 1037
rect 2830 861 2864 1037
rect 3012 861 3046 1037
rect 3130 861 3164 1037
rect 3312 861 3346 1037
rect 3430 861 3464 1037
rect 3612 861 3646 1037
rect 3730 861 3764 1037
rect 3912 861 3946 1037
rect 4030 861 4064 1037
rect 4212 861 4246 1037
rect 4330 861 4364 1037
rect 4512 861 4546 1037
rect 4630 861 4664 1037
rect 4812 861 4846 1037
rect 4930 861 4964 1037
rect 5112 861 5146 1037
rect 5230 861 5264 1037
rect 5412 861 5446 1037
rect 5530 861 5564 1037
rect 5712 861 5746 1037
rect 5830 861 5864 1037
rect 6012 861 6046 1037
rect 6130 861 6164 1037
rect 6312 861 6346 1037
rect 6430 861 6464 1037
rect 6612 861 6646 1037
rect 6730 861 6764 1037
rect 6912 861 6946 1037
rect 7030 861 7064 1037
rect 7212 861 7246 1037
rect 7330 861 7364 1037
rect 7512 861 7546 1037
rect 7630 861 7664 1037
rect 7812 861 7846 1037
rect 7930 861 7964 1037
rect 8112 861 8146 1037
rect 8230 861 8264 1037
rect 8412 861 8446 1037
rect 8530 861 8564 1037
rect 8712 861 8746 1037
rect 8830 861 8864 1037
rect 9012 861 9046 1037
rect 9130 861 9164 1037
rect 9312 861 9346 1037
rect 9430 861 9464 1037
rect 9612 861 9646 1037
rect 9730 861 9764 1037
rect 9912 861 9946 1037
rect 10030 861 10064 1037
rect 10212 861 10246 1037
rect 10330 861 10364 1037
rect 10512 861 10546 1037
rect 10630 861 10664 1037
rect 10812 861 10846 1037
rect 10930 861 10964 1037
rect 11112 861 11146 1037
rect 11230 861 11264 1037
rect 11412 861 11446 1037
rect 11530 861 11564 1037
rect 11712 861 11746 1037
rect 11830 861 11864 1037
rect 12012 861 12046 1037
rect 12130 861 12164 1037
rect 12312 861 12346 1037
rect 12430 861 12464 1037
rect 12612 861 12646 1037
rect 12730 861 12764 1037
rect 12912 861 12946 1037
rect 13030 861 13064 1037
rect 13212 861 13246 1037
rect 13330 861 13364 1037
rect 13512 861 13546 1037
rect 13630 861 13664 1037
rect 13812 861 13846 1037
rect 13930 861 13964 1037
rect 14112 861 14146 1037
rect 14230 861 14264 1037
rect 14412 861 14446 1037
rect 14530 861 14564 1037
rect 14712 861 14746 1037
rect 14830 861 14864 1037
rect 15012 861 15046 1037
rect 15130 861 15164 1037
rect 15312 861 15346 1037
<< mvpsubdiff >>
rect -14 508 15500 520
rect -14 474 124 508
rect 352 474 424 508
rect 652 474 724 508
rect 952 474 1024 508
rect 1252 474 1324 508
rect 1552 474 1624 508
rect 1852 474 1924 508
rect 2152 474 2224 508
rect 2452 474 2524 508
rect 2752 474 2824 508
rect 3052 474 3124 508
rect 3352 474 3424 508
rect 3652 474 3724 508
rect 3952 474 4024 508
rect 4252 474 4324 508
rect 4552 474 4624 508
rect 4852 474 4924 508
rect 5152 474 5224 508
rect 5452 474 5524 508
rect 5752 474 5824 508
rect 6052 474 6124 508
rect 6352 474 6424 508
rect 6652 474 6724 508
rect 6952 474 7024 508
rect 7252 474 7324 508
rect 7552 474 7624 508
rect 7852 474 7924 508
rect 8152 474 8224 508
rect 8452 474 8524 508
rect 8752 474 8824 508
rect 9052 474 9124 508
rect 9352 474 9424 508
rect 9652 474 9724 508
rect 9952 474 10024 508
rect 10252 474 10324 508
rect 10552 474 10624 508
rect 10852 474 10924 508
rect 11152 474 11224 508
rect 11452 474 11524 508
rect 11752 474 11824 508
rect 12052 474 12124 508
rect 12352 474 12424 508
rect 12652 474 12724 508
rect 12952 474 13024 508
rect 13252 474 13324 508
rect 13552 474 13624 508
rect 13852 474 13924 508
rect 14152 474 14224 508
rect 14452 474 14524 508
rect 14752 474 14824 508
rect 15052 474 15124 508
rect 15352 474 15500 508
rect -14 462 15500 474
rect -14 412 44 462
rect -14 144 -2 412
rect 32 144 44 412
rect 15442 412 15500 462
rect -14 94 44 144
rect 15442 144 15454 412
rect 15488 144 15500 412
rect 15442 94 15500 144
rect -14 82 15500 94
rect -14 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2524 82
rect 2752 48 2824 82
rect 3052 48 3124 82
rect 3352 48 3424 82
rect 3652 48 3724 82
rect 3952 48 4024 82
rect 4252 48 4324 82
rect 4552 48 4624 82
rect 4852 48 4924 82
rect 5152 48 5224 82
rect 5452 48 5524 82
rect 5752 48 5824 82
rect 6052 48 6124 82
rect 6352 48 6424 82
rect 6652 48 6724 82
rect 6952 48 7024 82
rect 7252 48 7324 82
rect 7552 48 7624 82
rect 7852 48 7924 82
rect 8152 48 8224 82
rect 8452 48 8524 82
rect 8752 48 8824 82
rect 9052 48 9124 82
rect 9352 48 9424 82
rect 9652 48 9724 82
rect 9952 48 10024 82
rect 10252 48 10324 82
rect 10552 48 10624 82
rect 10852 48 10924 82
rect 11152 48 11224 82
rect 11452 48 11524 82
rect 11752 48 11824 82
rect 12052 48 12124 82
rect 12352 48 12424 82
rect 12652 48 12724 82
rect 12952 48 13024 82
rect 13252 48 13324 82
rect 13552 48 13624 82
rect 13852 48 13924 82
rect 14152 48 14224 82
rect 14452 48 14524 82
rect 14752 48 14824 82
rect 15052 48 15124 82
rect 15352 48 15500 82
rect -14 36 15500 48
<< mvnsubdiff >>
rect 6 1214 15470 1226
rect 6 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2524 1214
rect 2752 1180 2824 1214
rect 3052 1180 3124 1214
rect 3352 1180 3424 1214
rect 3652 1180 3724 1214
rect 3952 1180 4024 1214
rect 4252 1180 4324 1214
rect 4552 1180 4624 1214
rect 4852 1180 4924 1214
rect 5152 1180 5224 1214
rect 5452 1180 5524 1214
rect 5752 1180 5824 1214
rect 6052 1180 6124 1214
rect 6352 1180 6424 1214
rect 6652 1180 6724 1214
rect 6952 1180 7024 1214
rect 7252 1180 7324 1214
rect 7552 1180 7624 1214
rect 7852 1180 7924 1214
rect 8152 1180 8224 1214
rect 8452 1180 8524 1214
rect 8752 1180 8824 1214
rect 9052 1180 9124 1214
rect 9352 1180 9424 1214
rect 9652 1180 9724 1214
rect 9952 1180 10024 1214
rect 10252 1180 10324 1214
rect 10552 1180 10624 1214
rect 10852 1180 10924 1214
rect 11152 1180 11224 1214
rect 11452 1180 11524 1214
rect 11752 1180 11824 1214
rect 12052 1180 12124 1214
rect 12352 1180 12424 1214
rect 12652 1180 12724 1214
rect 12952 1180 13024 1214
rect 13252 1180 13324 1214
rect 13552 1180 13624 1214
rect 13852 1180 13924 1214
rect 14152 1180 14224 1214
rect 14452 1180 14524 1214
rect 14752 1180 14824 1214
rect 15052 1180 15124 1214
rect 15352 1180 15470 1214
rect 6 1168 15470 1180
rect 6 1118 64 1168
rect 6 780 18 1118
rect 52 780 64 1118
rect 15412 1118 15470 1168
rect 6 730 64 780
rect 15412 780 15424 1118
rect 15458 780 15470 1118
rect 15412 730 15470 780
rect 6 718 15470 730
rect 6 684 124 718
rect 352 684 424 718
rect 652 684 724 718
rect 952 684 1024 718
rect 1252 684 1324 718
rect 1552 684 1624 718
rect 1852 684 1924 718
rect 2152 684 2224 718
rect 2452 684 2524 718
rect 2752 684 2824 718
rect 3052 684 3124 718
rect 3352 684 3424 718
rect 3652 684 3724 718
rect 3952 684 4024 718
rect 4252 684 4324 718
rect 4552 684 4624 718
rect 4852 684 4924 718
rect 5152 684 5224 718
rect 5452 684 5524 718
rect 5752 684 5824 718
rect 6052 684 6124 718
rect 6352 684 6424 718
rect 6652 684 6724 718
rect 6952 684 7024 718
rect 7252 684 7324 718
rect 7552 684 7624 718
rect 7852 684 7924 718
rect 8152 684 8224 718
rect 8452 684 8524 718
rect 8752 684 8824 718
rect 9052 684 9124 718
rect 9352 684 9424 718
rect 9652 684 9724 718
rect 9952 684 10024 718
rect 10252 684 10324 718
rect 10552 684 10624 718
rect 10852 684 10924 718
rect 11152 684 11224 718
rect 11452 684 11524 718
rect 11752 684 11824 718
rect 12052 684 12124 718
rect 12352 684 12424 718
rect 12652 684 12724 718
rect 12952 684 13024 718
rect 13252 684 13324 718
rect 13552 684 13624 718
rect 13852 684 13924 718
rect 14152 684 14224 718
rect 14452 684 14524 718
rect 14752 684 14824 718
rect 15052 684 15124 718
rect 15352 684 15470 718
rect 6 672 15470 684
<< mvpsubdiffcont >>
rect 124 474 352 508
rect 424 474 652 508
rect 724 474 952 508
rect 1024 474 1252 508
rect 1324 474 1552 508
rect 1624 474 1852 508
rect 1924 474 2152 508
rect 2224 474 2452 508
rect 2524 474 2752 508
rect 2824 474 3052 508
rect 3124 474 3352 508
rect 3424 474 3652 508
rect 3724 474 3952 508
rect 4024 474 4252 508
rect 4324 474 4552 508
rect 4624 474 4852 508
rect 4924 474 5152 508
rect 5224 474 5452 508
rect 5524 474 5752 508
rect 5824 474 6052 508
rect 6124 474 6352 508
rect 6424 474 6652 508
rect 6724 474 6952 508
rect 7024 474 7252 508
rect 7324 474 7552 508
rect 7624 474 7852 508
rect 7924 474 8152 508
rect 8224 474 8452 508
rect 8524 474 8752 508
rect 8824 474 9052 508
rect 9124 474 9352 508
rect 9424 474 9652 508
rect 9724 474 9952 508
rect 10024 474 10252 508
rect 10324 474 10552 508
rect 10624 474 10852 508
rect 10924 474 11152 508
rect 11224 474 11452 508
rect 11524 474 11752 508
rect 11824 474 12052 508
rect 12124 474 12352 508
rect 12424 474 12652 508
rect 12724 474 12952 508
rect 13024 474 13252 508
rect 13324 474 13552 508
rect 13624 474 13852 508
rect 13924 474 14152 508
rect 14224 474 14452 508
rect 14524 474 14752 508
rect 14824 474 15052 508
rect 15124 474 15352 508
rect -2 144 32 412
rect 15454 144 15488 412
rect 124 48 352 82
rect 424 48 652 82
rect 724 48 952 82
rect 1024 48 1252 82
rect 1324 48 1552 82
rect 1624 48 1852 82
rect 1924 48 2152 82
rect 2224 48 2452 82
rect 2524 48 2752 82
rect 2824 48 3052 82
rect 3124 48 3352 82
rect 3424 48 3652 82
rect 3724 48 3952 82
rect 4024 48 4252 82
rect 4324 48 4552 82
rect 4624 48 4852 82
rect 4924 48 5152 82
rect 5224 48 5452 82
rect 5524 48 5752 82
rect 5824 48 6052 82
rect 6124 48 6352 82
rect 6424 48 6652 82
rect 6724 48 6952 82
rect 7024 48 7252 82
rect 7324 48 7552 82
rect 7624 48 7852 82
rect 7924 48 8152 82
rect 8224 48 8452 82
rect 8524 48 8752 82
rect 8824 48 9052 82
rect 9124 48 9352 82
rect 9424 48 9652 82
rect 9724 48 9952 82
rect 10024 48 10252 82
rect 10324 48 10552 82
rect 10624 48 10852 82
rect 10924 48 11152 82
rect 11224 48 11452 82
rect 11524 48 11752 82
rect 11824 48 12052 82
rect 12124 48 12352 82
rect 12424 48 12652 82
rect 12724 48 12952 82
rect 13024 48 13252 82
rect 13324 48 13552 82
rect 13624 48 13852 82
rect 13924 48 14152 82
rect 14224 48 14452 82
rect 14524 48 14752 82
rect 14824 48 15052 82
rect 15124 48 15352 82
<< mvnsubdiffcont >>
rect 124 1180 352 1214
rect 424 1180 652 1214
rect 724 1180 952 1214
rect 1024 1180 1252 1214
rect 1324 1180 1552 1214
rect 1624 1180 1852 1214
rect 1924 1180 2152 1214
rect 2224 1180 2452 1214
rect 2524 1180 2752 1214
rect 2824 1180 3052 1214
rect 3124 1180 3352 1214
rect 3424 1180 3652 1214
rect 3724 1180 3952 1214
rect 4024 1180 4252 1214
rect 4324 1180 4552 1214
rect 4624 1180 4852 1214
rect 4924 1180 5152 1214
rect 5224 1180 5452 1214
rect 5524 1180 5752 1214
rect 5824 1180 6052 1214
rect 6124 1180 6352 1214
rect 6424 1180 6652 1214
rect 6724 1180 6952 1214
rect 7024 1180 7252 1214
rect 7324 1180 7552 1214
rect 7624 1180 7852 1214
rect 7924 1180 8152 1214
rect 8224 1180 8452 1214
rect 8524 1180 8752 1214
rect 8824 1180 9052 1214
rect 9124 1180 9352 1214
rect 9424 1180 9652 1214
rect 9724 1180 9952 1214
rect 10024 1180 10252 1214
rect 10324 1180 10552 1214
rect 10624 1180 10852 1214
rect 10924 1180 11152 1214
rect 11224 1180 11452 1214
rect 11524 1180 11752 1214
rect 11824 1180 12052 1214
rect 12124 1180 12352 1214
rect 12424 1180 12652 1214
rect 12724 1180 12952 1214
rect 13024 1180 13252 1214
rect 13324 1180 13552 1214
rect 13624 1180 13852 1214
rect 13924 1180 14152 1214
rect 14224 1180 14452 1214
rect 14524 1180 14752 1214
rect 14824 1180 15052 1214
rect 15124 1180 15352 1214
rect 18 780 52 1118
rect 15424 780 15458 1118
rect 124 684 352 718
rect 424 684 652 718
rect 724 684 952 718
rect 1024 684 1252 718
rect 1324 684 1552 718
rect 1624 684 1852 718
rect 1924 684 2152 718
rect 2224 684 2452 718
rect 2524 684 2752 718
rect 2824 684 3052 718
rect 3124 684 3352 718
rect 3424 684 3652 718
rect 3724 684 3952 718
rect 4024 684 4252 718
rect 4324 684 4552 718
rect 4624 684 4852 718
rect 4924 684 5152 718
rect 5224 684 5452 718
rect 5524 684 5752 718
rect 5824 684 6052 718
rect 6124 684 6352 718
rect 6424 684 6652 718
rect 6724 684 6952 718
rect 7024 684 7252 718
rect 7324 684 7552 718
rect 7624 684 7852 718
rect 7924 684 8152 718
rect 8224 684 8452 718
rect 8524 684 8752 718
rect 8824 684 9052 718
rect 9124 684 9352 718
rect 9424 684 9652 718
rect 9724 684 9952 718
rect 10024 684 10252 718
rect 10324 684 10552 718
rect 10624 684 10852 718
rect 10924 684 11152 718
rect 11224 684 11452 718
rect 11524 684 11752 718
rect 11824 684 12052 718
rect 12124 684 12352 718
rect 12424 684 12652 718
rect 12724 684 12952 718
rect 13024 684 13252 718
rect 13324 684 13552 718
rect 13624 684 13852 718
rect 13924 684 14152 718
rect 14224 684 14452 718
rect 14524 684 14752 718
rect 14824 684 15052 718
rect 15124 684 15352 718
<< poly >>
rect 188 1130 288 1146
rect 188 1096 204 1130
rect 272 1096 288 1130
rect 188 1049 288 1096
rect 488 1130 588 1146
rect 488 1096 504 1130
rect 572 1096 588 1130
rect 488 1049 588 1096
rect 788 1130 888 1146
rect 788 1096 804 1130
rect 872 1096 888 1130
rect 788 1049 888 1096
rect 1088 1130 1188 1146
rect 1088 1096 1104 1130
rect 1172 1096 1188 1130
rect 1088 1049 1188 1096
rect 1388 1130 1488 1146
rect 1388 1096 1404 1130
rect 1472 1096 1488 1130
rect 1388 1049 1488 1096
rect 1688 1130 1788 1146
rect 1688 1096 1704 1130
rect 1772 1096 1788 1130
rect 1688 1049 1788 1096
rect 1988 1130 2088 1146
rect 1988 1096 2004 1130
rect 2072 1096 2088 1130
rect 1988 1049 2088 1096
rect 2288 1130 2388 1146
rect 2288 1096 2304 1130
rect 2372 1096 2388 1130
rect 2288 1049 2388 1096
rect 2588 1130 2688 1146
rect 2588 1096 2604 1130
rect 2672 1096 2688 1130
rect 2588 1049 2688 1096
rect 2888 1130 2988 1146
rect 2888 1096 2904 1130
rect 2972 1096 2988 1130
rect 2888 1049 2988 1096
rect 3188 1130 3288 1146
rect 3188 1096 3204 1130
rect 3272 1096 3288 1130
rect 3188 1049 3288 1096
rect 3488 1130 3588 1146
rect 3488 1096 3504 1130
rect 3572 1096 3588 1130
rect 3488 1049 3588 1096
rect 3788 1130 3888 1146
rect 3788 1096 3804 1130
rect 3872 1096 3888 1130
rect 3788 1049 3888 1096
rect 4088 1130 4188 1146
rect 4088 1096 4104 1130
rect 4172 1096 4188 1130
rect 4088 1049 4188 1096
rect 4388 1130 4488 1146
rect 4388 1096 4404 1130
rect 4472 1096 4488 1130
rect 4388 1049 4488 1096
rect 4688 1130 4788 1146
rect 4688 1096 4704 1130
rect 4772 1096 4788 1130
rect 4688 1049 4788 1096
rect 4988 1130 5088 1146
rect 4988 1096 5004 1130
rect 5072 1096 5088 1130
rect 4988 1049 5088 1096
rect 5288 1130 5388 1146
rect 5288 1096 5304 1130
rect 5372 1096 5388 1130
rect 5288 1049 5388 1096
rect 5588 1130 5688 1146
rect 5588 1096 5604 1130
rect 5672 1096 5688 1130
rect 5588 1049 5688 1096
rect 5888 1130 5988 1146
rect 5888 1096 5904 1130
rect 5972 1096 5988 1130
rect 5888 1049 5988 1096
rect 6188 1130 6288 1146
rect 6188 1096 6204 1130
rect 6272 1096 6288 1130
rect 6188 1049 6288 1096
rect 6488 1130 6588 1146
rect 6488 1096 6504 1130
rect 6572 1096 6588 1130
rect 6488 1049 6588 1096
rect 6788 1130 6888 1146
rect 6788 1096 6804 1130
rect 6872 1096 6888 1130
rect 6788 1049 6888 1096
rect 7088 1130 7188 1146
rect 7088 1096 7104 1130
rect 7172 1096 7188 1130
rect 7088 1049 7188 1096
rect 7388 1130 7488 1146
rect 7388 1096 7404 1130
rect 7472 1096 7488 1130
rect 7388 1049 7488 1096
rect 7688 1130 7788 1146
rect 7688 1096 7704 1130
rect 7772 1096 7788 1130
rect 7688 1049 7788 1096
rect 7988 1130 8088 1146
rect 7988 1096 8004 1130
rect 8072 1096 8088 1130
rect 7988 1049 8088 1096
rect 8288 1130 8388 1146
rect 8288 1096 8304 1130
rect 8372 1096 8388 1130
rect 8288 1049 8388 1096
rect 8588 1130 8688 1146
rect 8588 1096 8604 1130
rect 8672 1096 8688 1130
rect 8588 1049 8688 1096
rect 8888 1130 8988 1146
rect 8888 1096 8904 1130
rect 8972 1096 8988 1130
rect 8888 1049 8988 1096
rect 9188 1130 9288 1146
rect 9188 1096 9204 1130
rect 9272 1096 9288 1130
rect 9188 1049 9288 1096
rect 9488 1130 9588 1146
rect 9488 1096 9504 1130
rect 9572 1096 9588 1130
rect 9488 1049 9588 1096
rect 9788 1130 9888 1146
rect 9788 1096 9804 1130
rect 9872 1096 9888 1130
rect 9788 1049 9888 1096
rect 10088 1130 10188 1146
rect 10088 1096 10104 1130
rect 10172 1096 10188 1130
rect 10088 1049 10188 1096
rect 10388 1130 10488 1146
rect 10388 1096 10404 1130
rect 10472 1096 10488 1130
rect 10388 1049 10488 1096
rect 10688 1130 10788 1146
rect 10688 1096 10704 1130
rect 10772 1096 10788 1130
rect 10688 1049 10788 1096
rect 10988 1130 11088 1146
rect 10988 1096 11004 1130
rect 11072 1096 11088 1130
rect 10988 1049 11088 1096
rect 11288 1130 11388 1146
rect 11288 1096 11304 1130
rect 11372 1096 11388 1130
rect 11288 1049 11388 1096
rect 11588 1130 11688 1146
rect 11588 1096 11604 1130
rect 11672 1096 11688 1130
rect 11588 1049 11688 1096
rect 11888 1130 11988 1146
rect 11888 1096 11904 1130
rect 11972 1096 11988 1130
rect 11888 1049 11988 1096
rect 12188 1130 12288 1146
rect 12188 1096 12204 1130
rect 12272 1096 12288 1130
rect 12188 1049 12288 1096
rect 12488 1130 12588 1146
rect 12488 1096 12504 1130
rect 12572 1096 12588 1130
rect 12488 1049 12588 1096
rect 12788 1130 12888 1146
rect 12788 1096 12804 1130
rect 12872 1096 12888 1130
rect 12788 1049 12888 1096
rect 13088 1130 13188 1146
rect 13088 1096 13104 1130
rect 13172 1096 13188 1130
rect 13088 1049 13188 1096
rect 13388 1130 13488 1146
rect 13388 1096 13404 1130
rect 13472 1096 13488 1130
rect 13388 1049 13488 1096
rect 13688 1130 13788 1146
rect 13688 1096 13704 1130
rect 13772 1096 13788 1130
rect 13688 1049 13788 1096
rect 13988 1130 14088 1146
rect 13988 1096 14004 1130
rect 14072 1096 14088 1130
rect 13988 1049 14088 1096
rect 14288 1130 14388 1146
rect 14288 1096 14304 1130
rect 14372 1096 14388 1130
rect 14288 1049 14388 1096
rect 14588 1130 14688 1146
rect 14588 1096 14604 1130
rect 14672 1096 14688 1130
rect 14588 1049 14688 1096
rect 14888 1130 14988 1146
rect 14888 1096 14904 1130
rect 14972 1096 14988 1130
rect 14888 1049 14988 1096
rect 15188 1130 15288 1146
rect 15188 1096 15204 1130
rect 15272 1096 15288 1130
rect 15188 1049 15288 1096
rect 188 802 288 849
rect 188 768 204 802
rect 272 768 288 802
rect 188 752 288 768
rect 488 802 588 849
rect 488 768 504 802
rect 572 768 588 802
rect 488 752 588 768
rect 788 802 888 849
rect 788 768 804 802
rect 872 768 888 802
rect 788 752 888 768
rect 1088 802 1188 849
rect 1088 768 1104 802
rect 1172 768 1188 802
rect 1088 752 1188 768
rect 1388 802 1488 849
rect 1388 768 1404 802
rect 1472 768 1488 802
rect 1388 752 1488 768
rect 1688 802 1788 849
rect 1688 768 1704 802
rect 1772 768 1788 802
rect 1688 752 1788 768
rect 1988 802 2088 849
rect 1988 768 2004 802
rect 2072 768 2088 802
rect 1988 752 2088 768
rect 2288 802 2388 849
rect 2288 768 2304 802
rect 2372 768 2388 802
rect 2288 752 2388 768
rect 2588 802 2688 849
rect 2588 768 2604 802
rect 2672 768 2688 802
rect 2588 752 2688 768
rect 2888 802 2988 849
rect 2888 768 2904 802
rect 2972 768 2988 802
rect 2888 752 2988 768
rect 3188 802 3288 849
rect 3188 768 3204 802
rect 3272 768 3288 802
rect 3188 752 3288 768
rect 3488 802 3588 849
rect 3488 768 3504 802
rect 3572 768 3588 802
rect 3488 752 3588 768
rect 3788 802 3888 849
rect 3788 768 3804 802
rect 3872 768 3888 802
rect 3788 752 3888 768
rect 4088 802 4188 849
rect 4088 768 4104 802
rect 4172 768 4188 802
rect 4088 752 4188 768
rect 4388 802 4488 849
rect 4388 768 4404 802
rect 4472 768 4488 802
rect 4388 752 4488 768
rect 4688 802 4788 849
rect 4688 768 4704 802
rect 4772 768 4788 802
rect 4688 752 4788 768
rect 4988 802 5088 849
rect 4988 768 5004 802
rect 5072 768 5088 802
rect 4988 752 5088 768
rect 5288 802 5388 849
rect 5288 768 5304 802
rect 5372 768 5388 802
rect 5288 752 5388 768
rect 5588 802 5688 849
rect 5588 768 5604 802
rect 5672 768 5688 802
rect 5588 752 5688 768
rect 5888 802 5988 849
rect 5888 768 5904 802
rect 5972 768 5988 802
rect 5888 752 5988 768
rect 6188 802 6288 849
rect 6188 768 6204 802
rect 6272 768 6288 802
rect 6188 752 6288 768
rect 6488 802 6588 849
rect 6488 768 6504 802
rect 6572 768 6588 802
rect 6488 752 6588 768
rect 6788 802 6888 849
rect 6788 768 6804 802
rect 6872 768 6888 802
rect 6788 752 6888 768
rect 7088 802 7188 849
rect 7088 768 7104 802
rect 7172 768 7188 802
rect 7088 752 7188 768
rect 7388 802 7488 849
rect 7388 768 7404 802
rect 7472 768 7488 802
rect 7388 752 7488 768
rect 7688 802 7788 849
rect 7688 768 7704 802
rect 7772 768 7788 802
rect 7688 752 7788 768
rect 7988 802 8088 849
rect 7988 768 8004 802
rect 8072 768 8088 802
rect 7988 752 8088 768
rect 8288 802 8388 849
rect 8288 768 8304 802
rect 8372 768 8388 802
rect 8288 752 8388 768
rect 8588 802 8688 849
rect 8588 768 8604 802
rect 8672 768 8688 802
rect 8588 752 8688 768
rect 8888 802 8988 849
rect 8888 768 8904 802
rect 8972 768 8988 802
rect 8888 752 8988 768
rect 9188 802 9288 849
rect 9188 768 9204 802
rect 9272 768 9288 802
rect 9188 752 9288 768
rect 9488 802 9588 849
rect 9488 768 9504 802
rect 9572 768 9588 802
rect 9488 752 9588 768
rect 9788 802 9888 849
rect 9788 768 9804 802
rect 9872 768 9888 802
rect 9788 752 9888 768
rect 10088 802 10188 849
rect 10088 768 10104 802
rect 10172 768 10188 802
rect 10088 752 10188 768
rect 10388 802 10488 849
rect 10388 768 10404 802
rect 10472 768 10488 802
rect 10388 752 10488 768
rect 10688 802 10788 849
rect 10688 768 10704 802
rect 10772 768 10788 802
rect 10688 752 10788 768
rect 10988 802 11088 849
rect 10988 768 11004 802
rect 11072 768 11088 802
rect 10988 752 11088 768
rect 11288 802 11388 849
rect 11288 768 11304 802
rect 11372 768 11388 802
rect 11288 752 11388 768
rect 11588 802 11688 849
rect 11588 768 11604 802
rect 11672 768 11688 802
rect 11588 752 11688 768
rect 11888 802 11988 849
rect 11888 768 11904 802
rect 11972 768 11988 802
rect 11888 752 11988 768
rect 12188 802 12288 849
rect 12188 768 12204 802
rect 12272 768 12288 802
rect 12188 752 12288 768
rect 12488 802 12588 849
rect 12488 768 12504 802
rect 12572 768 12588 802
rect 12488 752 12588 768
rect 12788 802 12888 849
rect 12788 768 12804 802
rect 12872 768 12888 802
rect 12788 752 12888 768
rect 13088 802 13188 849
rect 13088 768 13104 802
rect 13172 768 13188 802
rect 13088 752 13188 768
rect 13388 802 13488 849
rect 13388 768 13404 802
rect 13472 768 13488 802
rect 13388 752 13488 768
rect 13688 802 13788 849
rect 13688 768 13704 802
rect 13772 768 13788 802
rect 13688 752 13788 768
rect 13988 802 14088 849
rect 13988 768 14004 802
rect 14072 768 14088 802
rect 13988 752 14088 768
rect 14288 802 14388 849
rect 14288 768 14304 802
rect 14372 768 14388 802
rect 14288 752 14388 768
rect 14588 802 14688 849
rect 14588 768 14604 802
rect 14672 768 14688 802
rect 14588 752 14688 768
rect 14888 802 14988 849
rect 14888 768 14904 802
rect 14972 768 14988 802
rect 14888 752 14988 768
rect 15188 802 15288 849
rect 15188 768 15204 802
rect 15272 768 15288 802
rect 15188 752 15288 768
rect 188 415 288 431
rect 188 381 204 415
rect 272 381 288 415
rect 188 343 288 381
rect 488 415 588 431
rect 488 381 504 415
rect 572 381 588 415
rect 488 343 588 381
rect 788 415 888 431
rect 788 381 804 415
rect 872 381 888 415
rect 788 343 888 381
rect 1088 415 1188 431
rect 1088 381 1104 415
rect 1172 381 1188 415
rect 1088 343 1188 381
rect 1388 415 1488 431
rect 1388 381 1404 415
rect 1472 381 1488 415
rect 1388 343 1488 381
rect 1688 415 1788 431
rect 1688 381 1704 415
rect 1772 381 1788 415
rect 1688 343 1788 381
rect 1988 415 2088 431
rect 1988 381 2004 415
rect 2072 381 2088 415
rect 1988 343 2088 381
rect 2288 415 2388 431
rect 2288 381 2304 415
rect 2372 381 2388 415
rect 2288 343 2388 381
rect 2588 415 2688 431
rect 2588 381 2604 415
rect 2672 381 2688 415
rect 2588 343 2688 381
rect 2888 415 2988 431
rect 2888 381 2904 415
rect 2972 381 2988 415
rect 2888 343 2988 381
rect 3188 415 3288 431
rect 3188 381 3204 415
rect 3272 381 3288 415
rect 3188 343 3288 381
rect 3488 415 3588 431
rect 3488 381 3504 415
rect 3572 381 3588 415
rect 3488 343 3588 381
rect 3788 415 3888 431
rect 3788 381 3804 415
rect 3872 381 3888 415
rect 3788 343 3888 381
rect 4088 415 4188 431
rect 4088 381 4104 415
rect 4172 381 4188 415
rect 4088 343 4188 381
rect 4388 415 4488 431
rect 4388 381 4404 415
rect 4472 381 4488 415
rect 4388 343 4488 381
rect 4688 415 4788 431
rect 4688 381 4704 415
rect 4772 381 4788 415
rect 4688 343 4788 381
rect 4988 415 5088 431
rect 4988 381 5004 415
rect 5072 381 5088 415
rect 4988 343 5088 381
rect 5288 415 5388 431
rect 5288 381 5304 415
rect 5372 381 5388 415
rect 5288 343 5388 381
rect 5588 415 5688 431
rect 5588 381 5604 415
rect 5672 381 5688 415
rect 5588 343 5688 381
rect 5888 415 5988 431
rect 5888 381 5904 415
rect 5972 381 5988 415
rect 5888 343 5988 381
rect 6188 415 6288 431
rect 6188 381 6204 415
rect 6272 381 6288 415
rect 6188 343 6288 381
rect 6488 415 6588 431
rect 6488 381 6504 415
rect 6572 381 6588 415
rect 6488 343 6588 381
rect 6788 415 6888 431
rect 6788 381 6804 415
rect 6872 381 6888 415
rect 6788 343 6888 381
rect 7088 415 7188 431
rect 7088 381 7104 415
rect 7172 381 7188 415
rect 7088 343 7188 381
rect 7388 415 7488 431
rect 7388 381 7404 415
rect 7472 381 7488 415
rect 7388 343 7488 381
rect 7688 415 7788 431
rect 7688 381 7704 415
rect 7772 381 7788 415
rect 7688 343 7788 381
rect 7988 415 8088 431
rect 7988 381 8004 415
rect 8072 381 8088 415
rect 7988 343 8088 381
rect 8288 415 8388 431
rect 8288 381 8304 415
rect 8372 381 8388 415
rect 8288 343 8388 381
rect 8588 415 8688 431
rect 8588 381 8604 415
rect 8672 381 8688 415
rect 8588 343 8688 381
rect 8888 415 8988 431
rect 8888 381 8904 415
rect 8972 381 8988 415
rect 8888 343 8988 381
rect 9188 415 9288 431
rect 9188 381 9204 415
rect 9272 381 9288 415
rect 9188 343 9288 381
rect 9488 415 9588 431
rect 9488 381 9504 415
rect 9572 381 9588 415
rect 9488 343 9588 381
rect 9788 415 9888 431
rect 9788 381 9804 415
rect 9872 381 9888 415
rect 9788 343 9888 381
rect 10088 415 10188 431
rect 10088 381 10104 415
rect 10172 381 10188 415
rect 10088 343 10188 381
rect 10388 415 10488 431
rect 10388 381 10404 415
rect 10472 381 10488 415
rect 10388 343 10488 381
rect 10688 415 10788 431
rect 10688 381 10704 415
rect 10772 381 10788 415
rect 10688 343 10788 381
rect 10988 415 11088 431
rect 10988 381 11004 415
rect 11072 381 11088 415
rect 10988 343 11088 381
rect 11288 415 11388 431
rect 11288 381 11304 415
rect 11372 381 11388 415
rect 11288 343 11388 381
rect 11588 415 11688 431
rect 11588 381 11604 415
rect 11672 381 11688 415
rect 11588 343 11688 381
rect 11888 415 11988 431
rect 11888 381 11904 415
rect 11972 381 11988 415
rect 11888 343 11988 381
rect 12188 415 12288 431
rect 12188 381 12204 415
rect 12272 381 12288 415
rect 12188 343 12288 381
rect 12488 415 12588 431
rect 12488 381 12504 415
rect 12572 381 12588 415
rect 12488 343 12588 381
rect 12788 415 12888 431
rect 12788 381 12804 415
rect 12872 381 12888 415
rect 12788 343 12888 381
rect 13088 415 13188 431
rect 13088 381 13104 415
rect 13172 381 13188 415
rect 13088 343 13188 381
rect 13388 415 13488 431
rect 13388 381 13404 415
rect 13472 381 13488 415
rect 13388 343 13488 381
rect 13688 415 13788 431
rect 13688 381 13704 415
rect 13772 381 13788 415
rect 13688 343 13788 381
rect 13988 415 14088 431
rect 13988 381 14004 415
rect 14072 381 14088 415
rect 13988 343 14088 381
rect 14288 415 14388 431
rect 14288 381 14304 415
rect 14372 381 14388 415
rect 14288 343 14388 381
rect 14588 415 14688 431
rect 14588 381 14604 415
rect 14672 381 14688 415
rect 14588 343 14688 381
rect 14888 415 14988 431
rect 14888 381 14904 415
rect 14972 381 14988 415
rect 14888 343 14988 381
rect 15188 415 15288 431
rect 15188 381 15204 415
rect 15272 381 15288 415
rect 15188 343 15288 381
rect 188 175 288 213
rect 188 141 204 175
rect 272 141 288 175
rect 188 125 288 141
rect 488 175 588 213
rect 488 141 504 175
rect 572 141 588 175
rect 488 125 588 141
rect 788 175 888 213
rect 788 141 804 175
rect 872 141 888 175
rect 788 125 888 141
rect 1088 175 1188 213
rect 1088 141 1104 175
rect 1172 141 1188 175
rect 1088 125 1188 141
rect 1388 175 1488 213
rect 1388 141 1404 175
rect 1472 141 1488 175
rect 1388 125 1488 141
rect 1688 175 1788 213
rect 1688 141 1704 175
rect 1772 141 1788 175
rect 1688 125 1788 141
rect 1988 175 2088 213
rect 1988 141 2004 175
rect 2072 141 2088 175
rect 1988 125 2088 141
rect 2288 175 2388 213
rect 2288 141 2304 175
rect 2372 141 2388 175
rect 2288 125 2388 141
rect 2588 175 2688 213
rect 2588 141 2604 175
rect 2672 141 2688 175
rect 2588 125 2688 141
rect 2888 175 2988 213
rect 2888 141 2904 175
rect 2972 141 2988 175
rect 2888 125 2988 141
rect 3188 175 3288 213
rect 3188 141 3204 175
rect 3272 141 3288 175
rect 3188 125 3288 141
rect 3488 175 3588 213
rect 3488 141 3504 175
rect 3572 141 3588 175
rect 3488 125 3588 141
rect 3788 175 3888 213
rect 3788 141 3804 175
rect 3872 141 3888 175
rect 3788 125 3888 141
rect 4088 175 4188 213
rect 4088 141 4104 175
rect 4172 141 4188 175
rect 4088 125 4188 141
rect 4388 175 4488 213
rect 4388 141 4404 175
rect 4472 141 4488 175
rect 4388 125 4488 141
rect 4688 175 4788 213
rect 4688 141 4704 175
rect 4772 141 4788 175
rect 4688 125 4788 141
rect 4988 175 5088 213
rect 4988 141 5004 175
rect 5072 141 5088 175
rect 4988 125 5088 141
rect 5288 175 5388 213
rect 5288 141 5304 175
rect 5372 141 5388 175
rect 5288 125 5388 141
rect 5588 175 5688 213
rect 5588 141 5604 175
rect 5672 141 5688 175
rect 5588 125 5688 141
rect 5888 175 5988 213
rect 5888 141 5904 175
rect 5972 141 5988 175
rect 5888 125 5988 141
rect 6188 175 6288 213
rect 6188 141 6204 175
rect 6272 141 6288 175
rect 6188 125 6288 141
rect 6488 175 6588 213
rect 6488 141 6504 175
rect 6572 141 6588 175
rect 6488 125 6588 141
rect 6788 175 6888 213
rect 6788 141 6804 175
rect 6872 141 6888 175
rect 6788 125 6888 141
rect 7088 175 7188 213
rect 7088 141 7104 175
rect 7172 141 7188 175
rect 7088 125 7188 141
rect 7388 175 7488 213
rect 7388 141 7404 175
rect 7472 141 7488 175
rect 7388 125 7488 141
rect 7688 175 7788 213
rect 7688 141 7704 175
rect 7772 141 7788 175
rect 7688 125 7788 141
rect 7988 175 8088 213
rect 7988 141 8004 175
rect 8072 141 8088 175
rect 7988 125 8088 141
rect 8288 175 8388 213
rect 8288 141 8304 175
rect 8372 141 8388 175
rect 8288 125 8388 141
rect 8588 175 8688 213
rect 8588 141 8604 175
rect 8672 141 8688 175
rect 8588 125 8688 141
rect 8888 175 8988 213
rect 8888 141 8904 175
rect 8972 141 8988 175
rect 8888 125 8988 141
rect 9188 175 9288 213
rect 9188 141 9204 175
rect 9272 141 9288 175
rect 9188 125 9288 141
rect 9488 175 9588 213
rect 9488 141 9504 175
rect 9572 141 9588 175
rect 9488 125 9588 141
rect 9788 175 9888 213
rect 9788 141 9804 175
rect 9872 141 9888 175
rect 9788 125 9888 141
rect 10088 175 10188 213
rect 10088 141 10104 175
rect 10172 141 10188 175
rect 10088 125 10188 141
rect 10388 175 10488 213
rect 10388 141 10404 175
rect 10472 141 10488 175
rect 10388 125 10488 141
rect 10688 175 10788 213
rect 10688 141 10704 175
rect 10772 141 10788 175
rect 10688 125 10788 141
rect 10988 175 11088 213
rect 10988 141 11004 175
rect 11072 141 11088 175
rect 10988 125 11088 141
rect 11288 175 11388 213
rect 11288 141 11304 175
rect 11372 141 11388 175
rect 11288 125 11388 141
rect 11588 175 11688 213
rect 11588 141 11604 175
rect 11672 141 11688 175
rect 11588 125 11688 141
rect 11888 175 11988 213
rect 11888 141 11904 175
rect 11972 141 11988 175
rect 11888 125 11988 141
rect 12188 175 12288 213
rect 12188 141 12204 175
rect 12272 141 12288 175
rect 12188 125 12288 141
rect 12488 175 12588 213
rect 12488 141 12504 175
rect 12572 141 12588 175
rect 12488 125 12588 141
rect 12788 175 12888 213
rect 12788 141 12804 175
rect 12872 141 12888 175
rect 12788 125 12888 141
rect 13088 175 13188 213
rect 13088 141 13104 175
rect 13172 141 13188 175
rect 13088 125 13188 141
rect 13388 175 13488 213
rect 13388 141 13404 175
rect 13472 141 13488 175
rect 13388 125 13488 141
rect 13688 175 13788 213
rect 13688 141 13704 175
rect 13772 141 13788 175
rect 13688 125 13788 141
rect 13988 175 14088 213
rect 13988 141 14004 175
rect 14072 141 14088 175
rect 13988 125 14088 141
rect 14288 175 14388 213
rect 14288 141 14304 175
rect 14372 141 14388 175
rect 14288 125 14388 141
rect 14588 175 14688 213
rect 14588 141 14604 175
rect 14672 141 14688 175
rect 14588 125 14688 141
rect 14888 175 14988 213
rect 14888 141 14904 175
rect 14972 141 14988 175
rect 14888 125 14988 141
rect 15188 175 15288 213
rect 15188 141 15204 175
rect 15272 141 15288 175
rect 15188 125 15288 141
<< polycont >>
rect 204 1096 272 1130
rect 504 1096 572 1130
rect 804 1096 872 1130
rect 1104 1096 1172 1130
rect 1404 1096 1472 1130
rect 1704 1096 1772 1130
rect 2004 1096 2072 1130
rect 2304 1096 2372 1130
rect 2604 1096 2672 1130
rect 2904 1096 2972 1130
rect 3204 1096 3272 1130
rect 3504 1096 3572 1130
rect 3804 1096 3872 1130
rect 4104 1096 4172 1130
rect 4404 1096 4472 1130
rect 4704 1096 4772 1130
rect 5004 1096 5072 1130
rect 5304 1096 5372 1130
rect 5604 1096 5672 1130
rect 5904 1096 5972 1130
rect 6204 1096 6272 1130
rect 6504 1096 6572 1130
rect 6804 1096 6872 1130
rect 7104 1096 7172 1130
rect 7404 1096 7472 1130
rect 7704 1096 7772 1130
rect 8004 1096 8072 1130
rect 8304 1096 8372 1130
rect 8604 1096 8672 1130
rect 8904 1096 8972 1130
rect 9204 1096 9272 1130
rect 9504 1096 9572 1130
rect 9804 1096 9872 1130
rect 10104 1096 10172 1130
rect 10404 1096 10472 1130
rect 10704 1096 10772 1130
rect 11004 1096 11072 1130
rect 11304 1096 11372 1130
rect 11604 1096 11672 1130
rect 11904 1096 11972 1130
rect 12204 1096 12272 1130
rect 12504 1096 12572 1130
rect 12804 1096 12872 1130
rect 13104 1096 13172 1130
rect 13404 1096 13472 1130
rect 13704 1096 13772 1130
rect 14004 1096 14072 1130
rect 14304 1096 14372 1130
rect 14604 1096 14672 1130
rect 14904 1096 14972 1130
rect 15204 1096 15272 1130
rect 204 768 272 802
rect 504 768 572 802
rect 804 768 872 802
rect 1104 768 1172 802
rect 1404 768 1472 802
rect 1704 768 1772 802
rect 2004 768 2072 802
rect 2304 768 2372 802
rect 2604 768 2672 802
rect 2904 768 2972 802
rect 3204 768 3272 802
rect 3504 768 3572 802
rect 3804 768 3872 802
rect 4104 768 4172 802
rect 4404 768 4472 802
rect 4704 768 4772 802
rect 5004 768 5072 802
rect 5304 768 5372 802
rect 5604 768 5672 802
rect 5904 768 5972 802
rect 6204 768 6272 802
rect 6504 768 6572 802
rect 6804 768 6872 802
rect 7104 768 7172 802
rect 7404 768 7472 802
rect 7704 768 7772 802
rect 8004 768 8072 802
rect 8304 768 8372 802
rect 8604 768 8672 802
rect 8904 768 8972 802
rect 9204 768 9272 802
rect 9504 768 9572 802
rect 9804 768 9872 802
rect 10104 768 10172 802
rect 10404 768 10472 802
rect 10704 768 10772 802
rect 11004 768 11072 802
rect 11304 768 11372 802
rect 11604 768 11672 802
rect 11904 768 11972 802
rect 12204 768 12272 802
rect 12504 768 12572 802
rect 12804 768 12872 802
rect 13104 768 13172 802
rect 13404 768 13472 802
rect 13704 768 13772 802
rect 14004 768 14072 802
rect 14304 768 14372 802
rect 14604 768 14672 802
rect 14904 768 14972 802
rect 15204 768 15272 802
rect 204 381 272 415
rect 504 381 572 415
rect 804 381 872 415
rect 1104 381 1172 415
rect 1404 381 1472 415
rect 1704 381 1772 415
rect 2004 381 2072 415
rect 2304 381 2372 415
rect 2604 381 2672 415
rect 2904 381 2972 415
rect 3204 381 3272 415
rect 3504 381 3572 415
rect 3804 381 3872 415
rect 4104 381 4172 415
rect 4404 381 4472 415
rect 4704 381 4772 415
rect 5004 381 5072 415
rect 5304 381 5372 415
rect 5604 381 5672 415
rect 5904 381 5972 415
rect 6204 381 6272 415
rect 6504 381 6572 415
rect 6804 381 6872 415
rect 7104 381 7172 415
rect 7404 381 7472 415
rect 7704 381 7772 415
rect 8004 381 8072 415
rect 8304 381 8372 415
rect 8604 381 8672 415
rect 8904 381 8972 415
rect 9204 381 9272 415
rect 9504 381 9572 415
rect 9804 381 9872 415
rect 10104 381 10172 415
rect 10404 381 10472 415
rect 10704 381 10772 415
rect 11004 381 11072 415
rect 11304 381 11372 415
rect 11604 381 11672 415
rect 11904 381 11972 415
rect 12204 381 12272 415
rect 12504 381 12572 415
rect 12804 381 12872 415
rect 13104 381 13172 415
rect 13404 381 13472 415
rect 13704 381 13772 415
rect 14004 381 14072 415
rect 14304 381 14372 415
rect 14604 381 14672 415
rect 14904 381 14972 415
rect 15204 381 15272 415
rect 204 141 272 175
rect 504 141 572 175
rect 804 141 872 175
rect 1104 141 1172 175
rect 1404 141 1472 175
rect 1704 141 1772 175
rect 2004 141 2072 175
rect 2304 141 2372 175
rect 2604 141 2672 175
rect 2904 141 2972 175
rect 3204 141 3272 175
rect 3504 141 3572 175
rect 3804 141 3872 175
rect 4104 141 4172 175
rect 4404 141 4472 175
rect 4704 141 4772 175
rect 5004 141 5072 175
rect 5304 141 5372 175
rect 5604 141 5672 175
rect 5904 141 5972 175
rect 6204 141 6272 175
rect 6504 141 6572 175
rect 6804 141 6872 175
rect 7104 141 7172 175
rect 7404 141 7472 175
rect 7704 141 7772 175
rect 8004 141 8072 175
rect 8304 141 8372 175
rect 8604 141 8672 175
rect 8904 141 8972 175
rect 9204 141 9272 175
rect 9504 141 9572 175
rect 9804 141 9872 175
rect 10104 141 10172 175
rect 10404 141 10472 175
rect 10704 141 10772 175
rect 11004 141 11072 175
rect 11304 141 11372 175
rect 11604 141 11672 175
rect 11904 141 11972 175
rect 12204 141 12272 175
rect 12504 141 12572 175
rect 12804 141 12872 175
rect 13104 141 13172 175
rect 13404 141 13472 175
rect 13704 141 13772 175
rect 14004 141 14072 175
rect 14304 141 14372 175
rect 14604 141 14672 175
rect 14904 141 14972 175
rect 15204 141 15272 175
<< locali >>
rect 18 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2524 1214
rect 2752 1180 2824 1214
rect 3052 1180 3124 1214
rect 3352 1180 3424 1214
rect 3652 1180 3724 1214
rect 3952 1180 4024 1214
rect 4252 1180 4324 1214
rect 4552 1180 4624 1214
rect 4852 1180 4924 1214
rect 5152 1180 5224 1214
rect 5452 1180 5524 1214
rect 5752 1180 5824 1214
rect 6052 1180 6124 1214
rect 6352 1180 6424 1214
rect 6652 1180 6724 1214
rect 6952 1180 7024 1214
rect 7252 1180 7324 1214
rect 7552 1180 7624 1214
rect 7852 1180 7924 1214
rect 8152 1180 8224 1214
rect 8452 1180 8524 1214
rect 8752 1180 8824 1214
rect 9052 1180 9124 1214
rect 9352 1180 9424 1214
rect 9652 1180 9724 1214
rect 9952 1180 10024 1214
rect 10252 1180 10324 1214
rect 10552 1180 10624 1214
rect 10852 1180 10924 1214
rect 11152 1180 11224 1214
rect 11452 1180 11524 1214
rect 11752 1180 11824 1214
rect 12052 1180 12124 1214
rect 12352 1180 12424 1214
rect 12652 1180 12724 1214
rect 12952 1180 13024 1214
rect 13252 1180 13324 1214
rect 13552 1180 13624 1214
rect 13852 1180 13924 1214
rect 14152 1180 14224 1214
rect 14452 1180 14524 1214
rect 14752 1180 14824 1214
rect 15052 1180 15124 1214
rect 15352 1180 15458 1214
rect 18 1118 52 1180
rect 188 1096 204 1130
rect 272 1096 288 1130
rect 488 1096 504 1130
rect 572 1096 588 1130
rect 788 1096 804 1130
rect 872 1096 888 1130
rect 1088 1096 1104 1130
rect 1172 1096 1188 1130
rect 1388 1096 1404 1130
rect 1472 1096 1488 1130
rect 1688 1096 1704 1130
rect 1772 1096 1788 1130
rect 1988 1096 2004 1130
rect 2072 1096 2088 1130
rect 2288 1096 2304 1130
rect 2372 1096 2388 1130
rect 2588 1096 2604 1130
rect 2672 1096 2688 1130
rect 2888 1096 2904 1130
rect 2972 1096 2988 1130
rect 3188 1096 3204 1130
rect 3272 1096 3288 1130
rect 3488 1096 3504 1130
rect 3572 1096 3588 1130
rect 3788 1096 3804 1130
rect 3872 1096 3888 1130
rect 4088 1096 4104 1130
rect 4172 1096 4188 1130
rect 4388 1096 4404 1130
rect 4472 1096 4488 1130
rect 4688 1096 4704 1130
rect 4772 1096 4788 1130
rect 4988 1096 5004 1130
rect 5072 1096 5088 1130
rect 5288 1096 5304 1130
rect 5372 1096 5388 1130
rect 5588 1096 5604 1130
rect 5672 1096 5688 1130
rect 5888 1096 5904 1130
rect 5972 1096 5988 1130
rect 6188 1096 6204 1130
rect 6272 1096 6288 1130
rect 6488 1096 6504 1130
rect 6572 1096 6588 1130
rect 6788 1096 6804 1130
rect 6872 1096 6888 1130
rect 7088 1096 7104 1130
rect 7172 1096 7188 1130
rect 7388 1096 7404 1130
rect 7472 1096 7488 1130
rect 7688 1096 7704 1130
rect 7772 1096 7788 1130
rect 7988 1096 8004 1130
rect 8072 1096 8088 1130
rect 8288 1096 8304 1130
rect 8372 1096 8388 1130
rect 8588 1096 8604 1130
rect 8672 1096 8688 1130
rect 8888 1096 8904 1130
rect 8972 1096 8988 1130
rect 9188 1096 9204 1130
rect 9272 1096 9288 1130
rect 9488 1096 9504 1130
rect 9572 1096 9588 1130
rect 9788 1096 9804 1130
rect 9872 1096 9888 1130
rect 10088 1096 10104 1130
rect 10172 1096 10188 1130
rect 10388 1096 10404 1130
rect 10472 1096 10488 1130
rect 10688 1096 10704 1130
rect 10772 1096 10788 1130
rect 10988 1096 11004 1130
rect 11072 1096 11088 1130
rect 11288 1096 11304 1130
rect 11372 1096 11388 1130
rect 11588 1096 11604 1130
rect 11672 1096 11688 1130
rect 11888 1096 11904 1130
rect 11972 1096 11988 1130
rect 12188 1096 12204 1130
rect 12272 1096 12288 1130
rect 12488 1096 12504 1130
rect 12572 1096 12588 1130
rect 12788 1096 12804 1130
rect 12872 1096 12888 1130
rect 13088 1096 13104 1130
rect 13172 1096 13188 1130
rect 13388 1096 13404 1130
rect 13472 1096 13488 1130
rect 13688 1096 13704 1130
rect 13772 1096 13788 1130
rect 13988 1096 14004 1130
rect 14072 1096 14088 1130
rect 14288 1096 14304 1130
rect 14372 1096 14388 1130
rect 14588 1096 14604 1130
rect 14672 1096 14688 1130
rect 14888 1096 14904 1130
rect 14972 1096 14988 1130
rect 15188 1096 15204 1130
rect 15272 1096 15288 1130
rect 15424 1118 15458 1180
rect 130 1037 164 1053
rect 130 845 164 861
rect 312 1037 346 1053
rect 312 845 346 861
rect 430 1037 464 1053
rect 430 845 464 861
rect 612 1037 646 1053
rect 612 845 646 861
rect 730 1037 764 1053
rect 730 845 764 861
rect 912 1037 946 1053
rect 912 845 946 861
rect 1030 1037 1064 1053
rect 1030 845 1064 861
rect 1212 1037 1246 1053
rect 1212 845 1246 861
rect 1330 1037 1364 1053
rect 1330 845 1364 861
rect 1512 1037 1546 1053
rect 1512 845 1546 861
rect 1630 1037 1664 1053
rect 1630 845 1664 861
rect 1812 1037 1846 1053
rect 1812 845 1846 861
rect 1930 1037 1964 1053
rect 1930 845 1964 861
rect 2112 1037 2146 1053
rect 2112 845 2146 861
rect 2230 1037 2264 1053
rect 2230 845 2264 861
rect 2412 1037 2446 1053
rect 2412 845 2446 861
rect 2530 1037 2564 1053
rect 2530 845 2564 861
rect 2712 1037 2746 1053
rect 2712 845 2746 861
rect 2830 1037 2864 1053
rect 2830 845 2864 861
rect 3012 1037 3046 1053
rect 3012 845 3046 861
rect 3130 1037 3164 1053
rect 3130 845 3164 861
rect 3312 1037 3346 1053
rect 3312 845 3346 861
rect 3430 1037 3464 1053
rect 3430 845 3464 861
rect 3612 1037 3646 1053
rect 3612 845 3646 861
rect 3730 1037 3764 1053
rect 3730 845 3764 861
rect 3912 1037 3946 1053
rect 3912 845 3946 861
rect 4030 1037 4064 1053
rect 4030 845 4064 861
rect 4212 1037 4246 1053
rect 4212 845 4246 861
rect 4330 1037 4364 1053
rect 4330 845 4364 861
rect 4512 1037 4546 1053
rect 4512 845 4546 861
rect 4630 1037 4664 1053
rect 4630 845 4664 861
rect 4812 1037 4846 1053
rect 4812 845 4846 861
rect 4930 1037 4964 1053
rect 4930 845 4964 861
rect 5112 1037 5146 1053
rect 5112 845 5146 861
rect 5230 1037 5264 1053
rect 5230 845 5264 861
rect 5412 1037 5446 1053
rect 5412 845 5446 861
rect 5530 1037 5564 1053
rect 5530 845 5564 861
rect 5712 1037 5746 1053
rect 5712 845 5746 861
rect 5830 1037 5864 1053
rect 5830 845 5864 861
rect 6012 1037 6046 1053
rect 6012 845 6046 861
rect 6130 1037 6164 1053
rect 6130 845 6164 861
rect 6312 1037 6346 1053
rect 6312 845 6346 861
rect 6430 1037 6464 1053
rect 6430 845 6464 861
rect 6612 1037 6646 1053
rect 6612 845 6646 861
rect 6730 1037 6764 1053
rect 6730 845 6764 861
rect 6912 1037 6946 1053
rect 6912 845 6946 861
rect 7030 1037 7064 1053
rect 7030 845 7064 861
rect 7212 1037 7246 1053
rect 7212 845 7246 861
rect 7330 1037 7364 1053
rect 7330 845 7364 861
rect 7512 1037 7546 1053
rect 7512 845 7546 861
rect 7630 1037 7664 1053
rect 7630 845 7664 861
rect 7812 1037 7846 1053
rect 7812 845 7846 861
rect 7930 1037 7964 1053
rect 7930 845 7964 861
rect 8112 1037 8146 1053
rect 8112 845 8146 861
rect 8230 1037 8264 1053
rect 8230 845 8264 861
rect 8412 1037 8446 1053
rect 8412 845 8446 861
rect 8530 1037 8564 1053
rect 8530 845 8564 861
rect 8712 1037 8746 1053
rect 8712 845 8746 861
rect 8830 1037 8864 1053
rect 8830 845 8864 861
rect 9012 1037 9046 1053
rect 9012 845 9046 861
rect 9130 1037 9164 1053
rect 9130 845 9164 861
rect 9312 1037 9346 1053
rect 9312 845 9346 861
rect 9430 1037 9464 1053
rect 9430 845 9464 861
rect 9612 1037 9646 1053
rect 9612 845 9646 861
rect 9730 1037 9764 1053
rect 9730 845 9764 861
rect 9912 1037 9946 1053
rect 9912 845 9946 861
rect 10030 1037 10064 1053
rect 10030 845 10064 861
rect 10212 1037 10246 1053
rect 10212 845 10246 861
rect 10330 1037 10364 1053
rect 10330 845 10364 861
rect 10512 1037 10546 1053
rect 10512 845 10546 861
rect 10630 1037 10664 1053
rect 10630 845 10664 861
rect 10812 1037 10846 1053
rect 10812 845 10846 861
rect 10930 1037 10964 1053
rect 10930 845 10964 861
rect 11112 1037 11146 1053
rect 11112 845 11146 861
rect 11230 1037 11264 1053
rect 11230 845 11264 861
rect 11412 1037 11446 1053
rect 11412 845 11446 861
rect 11530 1037 11564 1053
rect 11530 845 11564 861
rect 11712 1037 11746 1053
rect 11712 845 11746 861
rect 11830 1037 11864 1053
rect 11830 845 11864 861
rect 12012 1037 12046 1053
rect 12012 845 12046 861
rect 12130 1037 12164 1053
rect 12130 845 12164 861
rect 12312 1037 12346 1053
rect 12312 845 12346 861
rect 12430 1037 12464 1053
rect 12430 845 12464 861
rect 12612 1037 12646 1053
rect 12612 845 12646 861
rect 12730 1037 12764 1053
rect 12730 845 12764 861
rect 12912 1037 12946 1053
rect 12912 845 12946 861
rect 13030 1037 13064 1053
rect 13030 845 13064 861
rect 13212 1037 13246 1053
rect 13212 845 13246 861
rect 13330 1037 13364 1053
rect 13330 845 13364 861
rect 13512 1037 13546 1053
rect 13512 845 13546 861
rect 13630 1037 13664 1053
rect 13630 845 13664 861
rect 13812 1037 13846 1053
rect 13812 845 13846 861
rect 13930 1037 13964 1053
rect 13930 845 13964 861
rect 14112 1037 14146 1053
rect 14112 845 14146 861
rect 14230 1037 14264 1053
rect 14230 845 14264 861
rect 14412 1037 14446 1053
rect 14412 845 14446 861
rect 14530 1037 14564 1053
rect 14530 845 14564 861
rect 14712 1037 14746 1053
rect 14712 845 14746 861
rect 14830 1037 14864 1053
rect 14830 845 14864 861
rect 15012 1037 15046 1053
rect 15012 845 15046 861
rect 15130 1037 15164 1053
rect 15130 845 15164 861
rect 15312 1037 15346 1053
rect 15312 845 15346 861
rect 18 718 52 780
rect 188 768 204 802
rect 272 768 288 802
rect 488 768 504 802
rect 572 768 588 802
rect 788 768 804 802
rect 872 768 888 802
rect 1088 768 1104 802
rect 1172 768 1188 802
rect 1388 768 1404 802
rect 1472 768 1488 802
rect 1688 768 1704 802
rect 1772 768 1788 802
rect 1988 768 2004 802
rect 2072 768 2088 802
rect 2288 768 2304 802
rect 2372 768 2388 802
rect 2588 768 2604 802
rect 2672 768 2688 802
rect 2888 768 2904 802
rect 2972 768 2988 802
rect 3188 768 3204 802
rect 3272 768 3288 802
rect 3488 768 3504 802
rect 3572 768 3588 802
rect 3788 768 3804 802
rect 3872 768 3888 802
rect 4088 768 4104 802
rect 4172 768 4188 802
rect 4388 768 4404 802
rect 4472 768 4488 802
rect 4688 768 4704 802
rect 4772 768 4788 802
rect 4988 768 5004 802
rect 5072 768 5088 802
rect 5288 768 5304 802
rect 5372 768 5388 802
rect 5588 768 5604 802
rect 5672 768 5688 802
rect 5888 768 5904 802
rect 5972 768 5988 802
rect 6188 768 6204 802
rect 6272 768 6288 802
rect 6488 768 6504 802
rect 6572 768 6588 802
rect 6788 768 6804 802
rect 6872 768 6888 802
rect 7088 768 7104 802
rect 7172 768 7188 802
rect 7388 768 7404 802
rect 7472 768 7488 802
rect 7688 768 7704 802
rect 7772 768 7788 802
rect 7988 768 8004 802
rect 8072 768 8088 802
rect 8288 768 8304 802
rect 8372 768 8388 802
rect 8588 768 8604 802
rect 8672 768 8688 802
rect 8888 768 8904 802
rect 8972 768 8988 802
rect 9188 768 9204 802
rect 9272 768 9288 802
rect 9488 768 9504 802
rect 9572 768 9588 802
rect 9788 768 9804 802
rect 9872 768 9888 802
rect 10088 768 10104 802
rect 10172 768 10188 802
rect 10388 768 10404 802
rect 10472 768 10488 802
rect 10688 768 10704 802
rect 10772 768 10788 802
rect 10988 768 11004 802
rect 11072 768 11088 802
rect 11288 768 11304 802
rect 11372 768 11388 802
rect 11588 768 11604 802
rect 11672 768 11688 802
rect 11888 768 11904 802
rect 11972 768 11988 802
rect 12188 768 12204 802
rect 12272 768 12288 802
rect 12488 768 12504 802
rect 12572 768 12588 802
rect 12788 768 12804 802
rect 12872 768 12888 802
rect 13088 768 13104 802
rect 13172 768 13188 802
rect 13388 768 13404 802
rect 13472 768 13488 802
rect 13688 768 13704 802
rect 13772 768 13788 802
rect 13988 768 14004 802
rect 14072 768 14088 802
rect 14288 768 14304 802
rect 14372 768 14388 802
rect 14588 768 14604 802
rect 14672 768 14688 802
rect 14888 768 14904 802
rect 14972 768 14988 802
rect 15188 768 15204 802
rect 15272 768 15288 802
rect 15424 718 15458 780
rect 18 684 124 718
rect 352 684 424 718
rect 652 684 724 718
rect 952 684 1024 718
rect 1252 684 1324 718
rect 1552 684 1624 718
rect 1852 684 1924 718
rect 2152 684 2224 718
rect 2452 684 2524 718
rect 2752 684 2824 718
rect 3052 684 3124 718
rect 3352 684 3424 718
rect 3652 684 3724 718
rect 3952 684 4024 718
rect 4252 684 4324 718
rect 4552 684 4624 718
rect 4852 684 4924 718
rect 5152 684 5224 718
rect 5452 684 5524 718
rect 5752 684 5824 718
rect 6052 684 6124 718
rect 6352 684 6424 718
rect 6652 684 6724 718
rect 6952 684 7024 718
rect 7252 684 7324 718
rect 7552 684 7624 718
rect 7852 684 7924 718
rect 8152 684 8224 718
rect 8452 684 8524 718
rect 8752 684 8824 718
rect 9052 684 9124 718
rect 9352 684 9424 718
rect 9652 684 9724 718
rect 9952 684 10024 718
rect 10252 684 10324 718
rect 10552 684 10624 718
rect 10852 684 10924 718
rect 11152 684 11224 718
rect 11452 684 11524 718
rect 11752 684 11824 718
rect 12052 684 12124 718
rect 12352 684 12424 718
rect 12652 684 12724 718
rect 12952 684 13024 718
rect 13252 684 13324 718
rect 13552 684 13624 718
rect 13852 684 13924 718
rect 14152 684 14224 718
rect 14452 684 14524 718
rect 14752 684 14824 718
rect 15052 684 15124 718
rect 15352 684 15458 718
rect -2 474 124 508
rect 352 474 424 508
rect 652 474 724 508
rect 952 474 1024 508
rect 1252 474 1324 508
rect 1552 474 1624 508
rect 1852 474 1924 508
rect 2152 474 2224 508
rect 2452 474 2524 508
rect 2752 474 2824 508
rect 3052 474 3124 508
rect 3352 474 3424 508
rect 3652 474 3724 508
rect 3952 474 4024 508
rect 4252 474 4324 508
rect 4552 474 4624 508
rect 4852 474 4924 508
rect 5152 474 5224 508
rect 5452 474 5524 508
rect 5752 474 5824 508
rect 6052 474 6124 508
rect 6352 474 6424 508
rect 6652 474 6724 508
rect 6952 474 7024 508
rect 7252 474 7324 508
rect 7552 474 7624 508
rect 7852 474 7924 508
rect 8152 474 8224 508
rect 8452 474 8524 508
rect 8752 474 8824 508
rect 9052 474 9124 508
rect 9352 474 9424 508
rect 9652 474 9724 508
rect 9952 474 10024 508
rect 10252 474 10324 508
rect 10552 474 10624 508
rect 10852 474 10924 508
rect 11152 474 11224 508
rect 11452 474 11524 508
rect 11752 474 11824 508
rect 12052 474 12124 508
rect 12352 474 12424 508
rect 12652 474 12724 508
rect 12952 474 13024 508
rect 13252 474 13324 508
rect 13552 474 13624 508
rect 13852 474 13924 508
rect 14152 474 14224 508
rect 14452 474 14524 508
rect 14752 474 14824 508
rect 15052 474 15124 508
rect 15352 474 15488 508
rect -2 412 32 474
rect 188 381 204 415
rect 272 381 288 415
rect 488 381 504 415
rect 572 381 588 415
rect 788 381 804 415
rect 872 381 888 415
rect 1088 381 1104 415
rect 1172 381 1188 415
rect 1388 381 1404 415
rect 1472 381 1488 415
rect 1688 381 1704 415
rect 1772 381 1788 415
rect 1988 381 2004 415
rect 2072 381 2088 415
rect 2288 381 2304 415
rect 2372 381 2388 415
rect 2588 381 2604 415
rect 2672 381 2688 415
rect 2888 381 2904 415
rect 2972 381 2988 415
rect 3188 381 3204 415
rect 3272 381 3288 415
rect 3488 381 3504 415
rect 3572 381 3588 415
rect 3788 381 3804 415
rect 3872 381 3888 415
rect 4088 381 4104 415
rect 4172 381 4188 415
rect 4388 381 4404 415
rect 4472 381 4488 415
rect 4688 381 4704 415
rect 4772 381 4788 415
rect 4988 381 5004 415
rect 5072 381 5088 415
rect 5288 381 5304 415
rect 5372 381 5388 415
rect 5588 381 5604 415
rect 5672 381 5688 415
rect 5888 381 5904 415
rect 5972 381 5988 415
rect 6188 381 6204 415
rect 6272 381 6288 415
rect 6488 381 6504 415
rect 6572 381 6588 415
rect 6788 381 6804 415
rect 6872 381 6888 415
rect 7088 381 7104 415
rect 7172 381 7188 415
rect 7388 381 7404 415
rect 7472 381 7488 415
rect 7688 381 7704 415
rect 7772 381 7788 415
rect 7988 381 8004 415
rect 8072 381 8088 415
rect 8288 381 8304 415
rect 8372 381 8388 415
rect 8588 381 8604 415
rect 8672 381 8688 415
rect 8888 381 8904 415
rect 8972 381 8988 415
rect 9188 381 9204 415
rect 9272 381 9288 415
rect 9488 381 9504 415
rect 9572 381 9588 415
rect 9788 381 9804 415
rect 9872 381 9888 415
rect 10088 381 10104 415
rect 10172 381 10188 415
rect 10388 381 10404 415
rect 10472 381 10488 415
rect 10688 381 10704 415
rect 10772 381 10788 415
rect 10988 381 11004 415
rect 11072 381 11088 415
rect 11288 381 11304 415
rect 11372 381 11388 415
rect 11588 381 11604 415
rect 11672 381 11688 415
rect 11888 381 11904 415
rect 11972 381 11988 415
rect 12188 381 12204 415
rect 12272 381 12288 415
rect 12488 381 12504 415
rect 12572 381 12588 415
rect 12788 381 12804 415
rect 12872 381 12888 415
rect 13088 381 13104 415
rect 13172 381 13188 415
rect 13388 381 13404 415
rect 13472 381 13488 415
rect 13688 381 13704 415
rect 13772 381 13788 415
rect 13988 381 14004 415
rect 14072 381 14088 415
rect 14288 381 14304 415
rect 14372 381 14388 415
rect 14588 381 14604 415
rect 14672 381 14688 415
rect 14888 381 14904 415
rect 14972 381 14988 415
rect 15188 381 15204 415
rect 15272 381 15288 415
rect 15454 412 15488 474
rect 130 331 164 347
rect 130 209 164 225
rect 312 331 346 347
rect 312 209 346 225
rect 430 331 464 347
rect 430 209 464 225
rect 612 331 646 347
rect 612 209 646 225
rect 730 331 764 347
rect 730 209 764 225
rect 912 331 946 347
rect 912 209 946 225
rect 1030 331 1064 347
rect 1030 209 1064 225
rect 1212 331 1246 347
rect 1212 209 1246 225
rect 1330 331 1364 347
rect 1330 209 1364 225
rect 1512 331 1546 347
rect 1512 209 1546 225
rect 1630 331 1664 347
rect 1630 209 1664 225
rect 1812 331 1846 347
rect 1812 209 1846 225
rect 1930 331 1964 347
rect 1930 209 1964 225
rect 2112 331 2146 347
rect 2112 209 2146 225
rect 2230 331 2264 347
rect 2230 209 2264 225
rect 2412 331 2446 347
rect 2412 209 2446 225
rect 2530 331 2564 347
rect 2530 209 2564 225
rect 2712 331 2746 347
rect 2712 209 2746 225
rect 2830 331 2864 347
rect 2830 209 2864 225
rect 3012 331 3046 347
rect 3012 209 3046 225
rect 3130 331 3164 347
rect 3130 209 3164 225
rect 3312 331 3346 347
rect 3312 209 3346 225
rect 3430 331 3464 347
rect 3430 209 3464 225
rect 3612 331 3646 347
rect 3612 209 3646 225
rect 3730 331 3764 347
rect 3730 209 3764 225
rect 3912 331 3946 347
rect 3912 209 3946 225
rect 4030 331 4064 347
rect 4030 209 4064 225
rect 4212 331 4246 347
rect 4212 209 4246 225
rect 4330 331 4364 347
rect 4330 209 4364 225
rect 4512 331 4546 347
rect 4512 209 4546 225
rect 4630 331 4664 347
rect 4630 209 4664 225
rect 4812 331 4846 347
rect 4812 209 4846 225
rect 4930 331 4964 347
rect 4930 209 4964 225
rect 5112 331 5146 347
rect 5112 209 5146 225
rect 5230 331 5264 347
rect 5230 209 5264 225
rect 5412 331 5446 347
rect 5412 209 5446 225
rect 5530 331 5564 347
rect 5530 209 5564 225
rect 5712 331 5746 347
rect 5712 209 5746 225
rect 5830 331 5864 347
rect 5830 209 5864 225
rect 6012 331 6046 347
rect 6012 209 6046 225
rect 6130 331 6164 347
rect 6130 209 6164 225
rect 6312 331 6346 347
rect 6312 209 6346 225
rect 6430 331 6464 347
rect 6430 209 6464 225
rect 6612 331 6646 347
rect 6612 209 6646 225
rect 6730 331 6764 347
rect 6730 209 6764 225
rect 6912 331 6946 347
rect 6912 209 6946 225
rect 7030 331 7064 347
rect 7030 209 7064 225
rect 7212 331 7246 347
rect 7212 209 7246 225
rect 7330 331 7364 347
rect 7330 209 7364 225
rect 7512 331 7546 347
rect 7512 209 7546 225
rect 7630 331 7664 347
rect 7630 209 7664 225
rect 7812 331 7846 347
rect 7812 209 7846 225
rect 7930 331 7964 347
rect 7930 209 7964 225
rect 8112 331 8146 347
rect 8112 209 8146 225
rect 8230 331 8264 347
rect 8230 209 8264 225
rect 8412 331 8446 347
rect 8412 209 8446 225
rect 8530 331 8564 347
rect 8530 209 8564 225
rect 8712 331 8746 347
rect 8712 209 8746 225
rect 8830 331 8864 347
rect 8830 209 8864 225
rect 9012 331 9046 347
rect 9012 209 9046 225
rect 9130 331 9164 347
rect 9130 209 9164 225
rect 9312 331 9346 347
rect 9312 209 9346 225
rect 9430 331 9464 347
rect 9430 209 9464 225
rect 9612 331 9646 347
rect 9612 209 9646 225
rect 9730 331 9764 347
rect 9730 209 9764 225
rect 9912 331 9946 347
rect 9912 209 9946 225
rect 10030 331 10064 347
rect 10030 209 10064 225
rect 10212 331 10246 347
rect 10212 209 10246 225
rect 10330 331 10364 347
rect 10330 209 10364 225
rect 10512 331 10546 347
rect 10512 209 10546 225
rect 10630 331 10664 347
rect 10630 209 10664 225
rect 10812 331 10846 347
rect 10812 209 10846 225
rect 10930 331 10964 347
rect 10930 209 10964 225
rect 11112 331 11146 347
rect 11112 209 11146 225
rect 11230 331 11264 347
rect 11230 209 11264 225
rect 11412 331 11446 347
rect 11412 209 11446 225
rect 11530 331 11564 347
rect 11530 209 11564 225
rect 11712 331 11746 347
rect 11712 209 11746 225
rect 11830 331 11864 347
rect 11830 209 11864 225
rect 12012 331 12046 347
rect 12012 209 12046 225
rect 12130 331 12164 347
rect 12130 209 12164 225
rect 12312 331 12346 347
rect 12312 209 12346 225
rect 12430 331 12464 347
rect 12430 209 12464 225
rect 12612 331 12646 347
rect 12612 209 12646 225
rect 12730 331 12764 347
rect 12730 209 12764 225
rect 12912 331 12946 347
rect 12912 209 12946 225
rect 13030 331 13064 347
rect 13030 209 13064 225
rect 13212 331 13246 347
rect 13212 209 13246 225
rect 13330 331 13364 347
rect 13330 209 13364 225
rect 13512 331 13546 347
rect 13512 209 13546 225
rect 13630 331 13664 347
rect 13630 209 13664 225
rect 13812 331 13846 347
rect 13812 209 13846 225
rect 13930 331 13964 347
rect 13930 209 13964 225
rect 14112 331 14146 347
rect 14112 209 14146 225
rect 14230 331 14264 347
rect 14230 209 14264 225
rect 14412 331 14446 347
rect 14412 209 14446 225
rect 14530 331 14564 347
rect 14530 209 14564 225
rect 14712 331 14746 347
rect 14712 209 14746 225
rect 14830 331 14864 347
rect 14830 209 14864 225
rect 15012 331 15046 347
rect 15012 209 15046 225
rect 15130 331 15164 347
rect 15130 209 15164 225
rect 15312 331 15346 347
rect 15312 209 15346 225
rect -2 82 32 144
rect 188 141 204 175
rect 272 141 288 175
rect 488 141 504 175
rect 572 141 588 175
rect 788 141 804 175
rect 872 141 888 175
rect 1088 141 1104 175
rect 1172 141 1188 175
rect 1388 141 1404 175
rect 1472 141 1488 175
rect 1688 141 1704 175
rect 1772 141 1788 175
rect 1988 141 2004 175
rect 2072 141 2088 175
rect 2288 141 2304 175
rect 2372 141 2388 175
rect 2588 141 2604 175
rect 2672 141 2688 175
rect 2888 141 2904 175
rect 2972 141 2988 175
rect 3188 141 3204 175
rect 3272 141 3288 175
rect 3488 141 3504 175
rect 3572 141 3588 175
rect 3788 141 3804 175
rect 3872 141 3888 175
rect 4088 141 4104 175
rect 4172 141 4188 175
rect 4388 141 4404 175
rect 4472 141 4488 175
rect 4688 141 4704 175
rect 4772 141 4788 175
rect 4988 141 5004 175
rect 5072 141 5088 175
rect 5288 141 5304 175
rect 5372 141 5388 175
rect 5588 141 5604 175
rect 5672 141 5688 175
rect 5888 141 5904 175
rect 5972 141 5988 175
rect 6188 141 6204 175
rect 6272 141 6288 175
rect 6488 141 6504 175
rect 6572 141 6588 175
rect 6788 141 6804 175
rect 6872 141 6888 175
rect 7088 141 7104 175
rect 7172 141 7188 175
rect 7388 141 7404 175
rect 7472 141 7488 175
rect 7688 141 7704 175
rect 7772 141 7788 175
rect 7988 141 8004 175
rect 8072 141 8088 175
rect 8288 141 8304 175
rect 8372 141 8388 175
rect 8588 141 8604 175
rect 8672 141 8688 175
rect 8888 141 8904 175
rect 8972 141 8988 175
rect 9188 141 9204 175
rect 9272 141 9288 175
rect 9488 141 9504 175
rect 9572 141 9588 175
rect 9788 141 9804 175
rect 9872 141 9888 175
rect 10088 141 10104 175
rect 10172 141 10188 175
rect 10388 141 10404 175
rect 10472 141 10488 175
rect 10688 141 10704 175
rect 10772 141 10788 175
rect 10988 141 11004 175
rect 11072 141 11088 175
rect 11288 141 11304 175
rect 11372 141 11388 175
rect 11588 141 11604 175
rect 11672 141 11688 175
rect 11888 141 11904 175
rect 11972 141 11988 175
rect 12188 141 12204 175
rect 12272 141 12288 175
rect 12488 141 12504 175
rect 12572 141 12588 175
rect 12788 141 12804 175
rect 12872 141 12888 175
rect 13088 141 13104 175
rect 13172 141 13188 175
rect 13388 141 13404 175
rect 13472 141 13488 175
rect 13688 141 13704 175
rect 13772 141 13788 175
rect 13988 141 14004 175
rect 14072 141 14088 175
rect 14288 141 14304 175
rect 14372 141 14388 175
rect 14588 141 14604 175
rect 14672 141 14688 175
rect 14888 141 14904 175
rect 14972 141 14988 175
rect 15188 141 15204 175
rect 15272 141 15288 175
rect 15454 82 15488 144
rect -2 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2524 82
rect 2752 48 2824 82
rect 3052 48 3124 82
rect 3352 48 3424 82
rect 3652 48 3724 82
rect 3952 48 4024 82
rect 4252 48 4324 82
rect 4552 48 4624 82
rect 4852 48 4924 82
rect 5152 48 5224 82
rect 5452 48 5524 82
rect 5752 48 5824 82
rect 6052 48 6124 82
rect 6352 48 6424 82
rect 6652 48 6724 82
rect 6952 48 7024 82
rect 7252 48 7324 82
rect 7552 48 7624 82
rect 7852 48 7924 82
rect 8152 48 8224 82
rect 8452 48 8524 82
rect 8752 48 8824 82
rect 9052 48 9124 82
rect 9352 48 9424 82
rect 9652 48 9724 82
rect 9952 48 10024 82
rect 10252 48 10324 82
rect 10552 48 10624 82
rect 10852 48 10924 82
rect 11152 48 11224 82
rect 11452 48 11524 82
rect 11752 48 11824 82
rect 12052 48 12124 82
rect 12352 48 12424 82
rect 12652 48 12724 82
rect 12952 48 13024 82
rect 13252 48 13324 82
rect 13552 48 13624 82
rect 13852 48 13924 82
rect 14152 48 14224 82
rect 14452 48 14524 82
rect 14752 48 14824 82
rect 15052 48 15124 82
rect 15352 48 15488 82
<< viali >>
rect 124 1180 352 1214
rect 424 1180 652 1214
rect 724 1180 952 1214
rect 1024 1180 1252 1214
rect 1324 1180 1552 1214
rect 1624 1180 1852 1214
rect 1924 1180 2152 1214
rect 2224 1180 2452 1214
rect 2524 1180 2752 1214
rect 2824 1180 3052 1214
rect 3124 1180 3352 1214
rect 3424 1180 3652 1214
rect 3724 1180 3952 1214
rect 4024 1180 4252 1214
rect 4324 1180 4552 1214
rect 4624 1180 4852 1214
rect 4924 1180 5152 1214
rect 5224 1180 5452 1214
rect 5524 1180 5752 1214
rect 5824 1180 6052 1214
rect 6124 1180 6352 1214
rect 6424 1180 6652 1214
rect 6724 1180 6952 1214
rect 7024 1180 7252 1214
rect 7324 1180 7552 1214
rect 7624 1180 7852 1214
rect 7924 1180 8152 1214
rect 8224 1180 8452 1214
rect 8524 1180 8752 1214
rect 8824 1180 9052 1214
rect 9124 1180 9352 1214
rect 9424 1180 9652 1214
rect 9724 1180 9952 1214
rect 10024 1180 10252 1214
rect 10324 1180 10552 1214
rect 10624 1180 10852 1214
rect 10924 1180 11152 1214
rect 11224 1180 11452 1214
rect 11524 1180 11752 1214
rect 11824 1180 12052 1214
rect 12124 1180 12352 1214
rect 12424 1180 12652 1214
rect 12724 1180 12952 1214
rect 13024 1180 13252 1214
rect 13324 1180 13552 1214
rect 13624 1180 13852 1214
rect 13924 1180 14152 1214
rect 14224 1180 14452 1214
rect 14524 1180 14752 1214
rect 14824 1180 15052 1214
rect 15124 1180 15352 1214
rect 204 1096 272 1130
rect 504 1096 572 1130
rect 804 1096 872 1130
rect 1104 1096 1172 1130
rect 1404 1096 1472 1130
rect 1704 1096 1772 1130
rect 2004 1096 2072 1130
rect 2304 1096 2372 1130
rect 2604 1096 2672 1130
rect 2904 1096 2972 1130
rect 3204 1096 3272 1130
rect 3504 1096 3572 1130
rect 3804 1096 3872 1130
rect 4104 1096 4172 1130
rect 4404 1096 4472 1130
rect 4704 1096 4772 1130
rect 5004 1096 5072 1130
rect 5304 1096 5372 1130
rect 5604 1096 5672 1130
rect 5904 1096 5972 1130
rect 6204 1096 6272 1130
rect 6504 1096 6572 1130
rect 6804 1096 6872 1130
rect 7104 1096 7172 1130
rect 7404 1096 7472 1130
rect 7704 1096 7772 1130
rect 8004 1096 8072 1130
rect 8304 1096 8372 1130
rect 8604 1096 8672 1130
rect 8904 1096 8972 1130
rect 9204 1096 9272 1130
rect 9504 1096 9572 1130
rect 9804 1096 9872 1130
rect 10104 1096 10172 1130
rect 10404 1096 10472 1130
rect 10704 1096 10772 1130
rect 11004 1096 11072 1130
rect 11304 1096 11372 1130
rect 11604 1096 11672 1130
rect 11904 1096 11972 1130
rect 12204 1096 12272 1130
rect 12504 1096 12572 1130
rect 12804 1096 12872 1130
rect 13104 1096 13172 1130
rect 13404 1096 13472 1130
rect 13704 1096 13772 1130
rect 14004 1096 14072 1130
rect 14304 1096 14372 1130
rect 14604 1096 14672 1130
rect 14904 1096 14972 1130
rect 15204 1096 15272 1130
rect 130 861 164 1037
rect 312 861 346 1037
rect 430 861 464 1037
rect 612 861 646 1037
rect 730 861 764 1037
rect 912 861 946 1037
rect 1030 861 1064 1037
rect 1212 861 1246 1037
rect 1330 861 1364 1037
rect 1512 861 1546 1037
rect 1630 861 1664 1037
rect 1812 861 1846 1037
rect 1930 861 1964 1037
rect 2112 861 2146 1037
rect 2230 861 2264 1037
rect 2412 861 2446 1037
rect 2530 861 2564 1037
rect 2712 861 2746 1037
rect 2830 861 2864 1037
rect 3012 861 3046 1037
rect 3130 861 3164 1037
rect 3312 861 3346 1037
rect 3430 861 3464 1037
rect 3612 861 3646 1037
rect 3730 861 3764 1037
rect 3912 861 3946 1037
rect 4030 861 4064 1037
rect 4212 861 4246 1037
rect 4330 861 4364 1037
rect 4512 861 4546 1037
rect 4630 861 4664 1037
rect 4812 861 4846 1037
rect 4930 861 4964 1037
rect 5112 861 5146 1037
rect 5230 861 5264 1037
rect 5412 861 5446 1037
rect 5530 861 5564 1037
rect 5712 861 5746 1037
rect 5830 861 5864 1037
rect 6012 861 6046 1037
rect 6130 861 6164 1037
rect 6312 861 6346 1037
rect 6430 861 6464 1037
rect 6612 861 6646 1037
rect 6730 861 6764 1037
rect 6912 861 6946 1037
rect 7030 861 7064 1037
rect 7212 861 7246 1037
rect 7330 861 7364 1037
rect 7512 861 7546 1037
rect 7630 861 7664 1037
rect 7812 861 7846 1037
rect 7930 861 7964 1037
rect 8112 861 8146 1037
rect 8230 861 8264 1037
rect 8412 861 8446 1037
rect 8530 861 8564 1037
rect 8712 861 8746 1037
rect 8830 861 8864 1037
rect 9012 861 9046 1037
rect 9130 861 9164 1037
rect 9312 861 9346 1037
rect 9430 861 9464 1037
rect 9612 861 9646 1037
rect 9730 861 9764 1037
rect 9912 861 9946 1037
rect 10030 861 10064 1037
rect 10212 861 10246 1037
rect 10330 861 10364 1037
rect 10512 861 10546 1037
rect 10630 861 10664 1037
rect 10812 861 10846 1037
rect 10930 861 10964 1037
rect 11112 861 11146 1037
rect 11230 861 11264 1037
rect 11412 861 11446 1037
rect 11530 861 11564 1037
rect 11712 861 11746 1037
rect 11830 861 11864 1037
rect 12012 861 12046 1037
rect 12130 861 12164 1037
rect 12312 861 12346 1037
rect 12430 861 12464 1037
rect 12612 861 12646 1037
rect 12730 861 12764 1037
rect 12912 861 12946 1037
rect 13030 861 13064 1037
rect 13212 861 13246 1037
rect 13330 861 13364 1037
rect 13512 861 13546 1037
rect 13630 861 13664 1037
rect 13812 861 13846 1037
rect 13930 861 13964 1037
rect 14112 861 14146 1037
rect 14230 861 14264 1037
rect 14412 861 14446 1037
rect 14530 861 14564 1037
rect 14712 861 14746 1037
rect 14830 861 14864 1037
rect 15012 861 15046 1037
rect 15130 861 15164 1037
rect 15312 861 15346 1037
rect 204 768 272 802
rect 504 768 572 802
rect 804 768 872 802
rect 1104 768 1172 802
rect 1404 768 1472 802
rect 1704 768 1772 802
rect 2004 768 2072 802
rect 2304 768 2372 802
rect 2604 768 2672 802
rect 2904 768 2972 802
rect 3204 768 3272 802
rect 3504 768 3572 802
rect 3804 768 3872 802
rect 4104 768 4172 802
rect 4404 768 4472 802
rect 4704 768 4772 802
rect 5004 768 5072 802
rect 5304 768 5372 802
rect 5604 768 5672 802
rect 5904 768 5972 802
rect 6204 768 6272 802
rect 6504 768 6572 802
rect 6804 768 6872 802
rect 7104 768 7172 802
rect 7404 768 7472 802
rect 7704 768 7772 802
rect 8004 768 8072 802
rect 8304 768 8372 802
rect 8604 768 8672 802
rect 8904 768 8972 802
rect 9204 768 9272 802
rect 9504 768 9572 802
rect 9804 768 9872 802
rect 10104 768 10172 802
rect 10404 768 10472 802
rect 10704 768 10772 802
rect 11004 768 11072 802
rect 11304 768 11372 802
rect 11604 768 11672 802
rect 11904 768 11972 802
rect 12204 768 12272 802
rect 12504 768 12572 802
rect 12804 768 12872 802
rect 13104 768 13172 802
rect 13404 768 13472 802
rect 13704 768 13772 802
rect 14004 768 14072 802
rect 14304 768 14372 802
rect 14604 768 14672 802
rect 14904 768 14972 802
rect 15204 768 15272 802
rect 204 381 272 415
rect 504 381 572 415
rect 804 381 872 415
rect 1104 381 1172 415
rect 1404 381 1472 415
rect 1704 381 1772 415
rect 2004 381 2072 415
rect 2304 381 2372 415
rect 2604 381 2672 415
rect 2904 381 2972 415
rect 3204 381 3272 415
rect 3504 381 3572 415
rect 3804 381 3872 415
rect 4104 381 4172 415
rect 4404 381 4472 415
rect 4704 381 4772 415
rect 5004 381 5072 415
rect 5304 381 5372 415
rect 5604 381 5672 415
rect 5904 381 5972 415
rect 6204 381 6272 415
rect 6504 381 6572 415
rect 6804 381 6872 415
rect 7104 381 7172 415
rect 7404 381 7472 415
rect 7704 381 7772 415
rect 8004 381 8072 415
rect 8304 381 8372 415
rect 8604 381 8672 415
rect 8904 381 8972 415
rect 9204 381 9272 415
rect 9504 381 9572 415
rect 9804 381 9872 415
rect 10104 381 10172 415
rect 10404 381 10472 415
rect 10704 381 10772 415
rect 11004 381 11072 415
rect 11304 381 11372 415
rect 11604 381 11672 415
rect 11904 381 11972 415
rect 12204 381 12272 415
rect 12504 381 12572 415
rect 12804 381 12872 415
rect 13104 381 13172 415
rect 13404 381 13472 415
rect 13704 381 13772 415
rect 14004 381 14072 415
rect 14304 381 14372 415
rect 14604 381 14672 415
rect 14904 381 14972 415
rect 15204 381 15272 415
rect 130 225 164 331
rect 312 225 346 331
rect 430 225 464 331
rect 612 225 646 331
rect 730 225 764 331
rect 912 225 946 331
rect 1030 225 1064 331
rect 1212 225 1246 331
rect 1330 225 1364 331
rect 1512 225 1546 331
rect 1630 225 1664 331
rect 1812 225 1846 331
rect 1930 225 1964 331
rect 2112 225 2146 331
rect 2230 225 2264 331
rect 2412 225 2446 331
rect 2530 225 2564 331
rect 2712 225 2746 331
rect 2830 225 2864 331
rect 3012 225 3046 331
rect 3130 225 3164 331
rect 3312 225 3346 331
rect 3430 225 3464 331
rect 3612 225 3646 331
rect 3730 225 3764 331
rect 3912 225 3946 331
rect 4030 225 4064 331
rect 4212 225 4246 331
rect 4330 225 4364 331
rect 4512 225 4546 331
rect 4630 225 4664 331
rect 4812 225 4846 331
rect 4930 225 4964 331
rect 5112 225 5146 331
rect 5230 225 5264 331
rect 5412 225 5446 331
rect 5530 225 5564 331
rect 5712 225 5746 331
rect 5830 225 5864 331
rect 6012 225 6046 331
rect 6130 225 6164 331
rect 6312 225 6346 331
rect 6430 225 6464 331
rect 6612 225 6646 331
rect 6730 225 6764 331
rect 6912 225 6946 331
rect 7030 225 7064 331
rect 7212 225 7246 331
rect 7330 225 7364 331
rect 7512 225 7546 331
rect 7630 225 7664 331
rect 7812 225 7846 331
rect 7930 225 7964 331
rect 8112 225 8146 331
rect 8230 225 8264 331
rect 8412 225 8446 331
rect 8530 225 8564 331
rect 8712 225 8746 331
rect 8830 225 8864 331
rect 9012 225 9046 331
rect 9130 225 9164 331
rect 9312 225 9346 331
rect 9430 225 9464 331
rect 9612 225 9646 331
rect 9730 225 9764 331
rect 9912 225 9946 331
rect 10030 225 10064 331
rect 10212 225 10246 331
rect 10330 225 10364 331
rect 10512 225 10546 331
rect 10630 225 10664 331
rect 10812 225 10846 331
rect 10930 225 10964 331
rect 11112 225 11146 331
rect 11230 225 11264 331
rect 11412 225 11446 331
rect 11530 225 11564 331
rect 11712 225 11746 331
rect 11830 225 11864 331
rect 12012 225 12046 331
rect 12130 225 12164 331
rect 12312 225 12346 331
rect 12430 225 12464 331
rect 12612 225 12646 331
rect 12730 225 12764 331
rect 12912 225 12946 331
rect 13030 225 13064 331
rect 13212 225 13246 331
rect 13330 225 13364 331
rect 13512 225 13546 331
rect 13630 225 13664 331
rect 13812 225 13846 331
rect 13930 225 13964 331
rect 14112 225 14146 331
rect 14230 225 14264 331
rect 14412 225 14446 331
rect 14530 225 14564 331
rect 14712 225 14746 331
rect 14830 225 14864 331
rect 15012 225 15046 331
rect 15130 225 15164 331
rect 15312 225 15346 331
rect 204 141 272 175
rect 504 141 572 175
rect 804 141 872 175
rect 1104 141 1172 175
rect 1404 141 1472 175
rect 1704 141 1772 175
rect 2004 141 2072 175
rect 2304 141 2372 175
rect 2604 141 2672 175
rect 2904 141 2972 175
rect 3204 141 3272 175
rect 3504 141 3572 175
rect 3804 141 3872 175
rect 4104 141 4172 175
rect 4404 141 4472 175
rect 4704 141 4772 175
rect 5004 141 5072 175
rect 5304 141 5372 175
rect 5604 141 5672 175
rect 5904 141 5972 175
rect 6204 141 6272 175
rect 6504 141 6572 175
rect 6804 141 6872 175
rect 7104 141 7172 175
rect 7404 141 7472 175
rect 7704 141 7772 175
rect 8004 141 8072 175
rect 8304 141 8372 175
rect 8604 141 8672 175
rect 8904 141 8972 175
rect 9204 141 9272 175
rect 9504 141 9572 175
rect 9804 141 9872 175
rect 10104 141 10172 175
rect 10404 141 10472 175
rect 10704 141 10772 175
rect 11004 141 11072 175
rect 11304 141 11372 175
rect 11604 141 11672 175
rect 11904 141 11972 175
rect 12204 141 12272 175
rect 12504 141 12572 175
rect 12804 141 12872 175
rect 13104 141 13172 175
rect 13404 141 13472 175
rect 13704 141 13772 175
rect 14004 141 14072 175
rect 14304 141 14372 175
rect 14604 141 14672 175
rect 14904 141 14972 175
rect 15204 141 15272 175
rect 124 48 352 82
rect 424 48 652 82
rect 724 48 952 82
rect 1024 48 1252 82
rect 1324 48 1552 82
rect 1624 48 1852 82
rect 1924 48 2152 82
rect 2224 48 2452 82
rect 2524 48 2752 82
rect 2824 48 3052 82
rect 3124 48 3352 82
rect 3424 48 3652 82
rect 3724 48 3952 82
rect 4024 48 4252 82
rect 4324 48 4552 82
rect 4624 48 4852 82
rect 4924 48 5152 82
rect 5224 48 5452 82
rect 5524 48 5752 82
rect 5824 48 6052 82
rect 6124 48 6352 82
rect 6424 48 6652 82
rect 6724 48 6952 82
rect 7024 48 7252 82
rect 7324 48 7552 82
rect 7624 48 7852 82
rect 7924 48 8152 82
rect 8224 48 8452 82
rect 8524 48 8752 82
rect 8824 48 9052 82
rect 9124 48 9352 82
rect 9424 48 9652 82
rect 9724 48 9952 82
rect 10024 48 10252 82
rect 10324 48 10552 82
rect 10624 48 10852 82
rect 10924 48 11152 82
rect 11224 48 11452 82
rect 11524 48 11752 82
rect 11824 48 12052 82
rect 12124 48 12352 82
rect 12424 48 12652 82
rect 12724 48 12952 82
rect 13024 48 13252 82
rect 13324 48 13552 82
rect 13624 48 13852 82
rect 13924 48 14152 82
rect 14224 48 14452 82
rect 14524 48 14752 82
rect 14824 48 15052 82
rect 15124 48 15352 82
<< metal1 >>
rect 88 1214 15388 1226
rect 88 1180 124 1214
rect 352 1180 424 1214
rect 652 1180 724 1214
rect 952 1180 1024 1214
rect 1252 1180 1324 1214
rect 1552 1180 1624 1214
rect 1852 1180 1924 1214
rect 2152 1180 2224 1214
rect 2452 1180 2524 1214
rect 2752 1180 2824 1214
rect 3052 1180 3124 1214
rect 3352 1180 3424 1214
rect 3652 1180 3724 1214
rect 3952 1180 4024 1214
rect 4252 1180 4324 1214
rect 4552 1180 4624 1214
rect 4852 1180 4924 1214
rect 5152 1180 5224 1214
rect 5452 1180 5524 1214
rect 5752 1180 5824 1214
rect 6052 1180 6124 1214
rect 6352 1180 6424 1214
rect 6652 1180 6724 1214
rect 6952 1180 7024 1214
rect 7252 1180 7324 1214
rect 7552 1180 7624 1214
rect 7852 1180 7924 1214
rect 8152 1180 8224 1214
rect 8452 1180 8524 1214
rect 8752 1180 8824 1214
rect 9052 1180 9124 1214
rect 9352 1180 9424 1214
rect 9652 1180 9724 1214
rect 9952 1180 10024 1214
rect 10252 1180 10324 1214
rect 10552 1180 10624 1214
rect 10852 1180 10924 1214
rect 11152 1180 11224 1214
rect 11452 1180 11524 1214
rect 11752 1180 11824 1214
rect 12052 1180 12124 1214
rect 12352 1180 12424 1214
rect 12652 1180 12724 1214
rect 12952 1180 13024 1214
rect 13252 1180 13324 1214
rect 13552 1180 13624 1214
rect 13852 1180 13924 1214
rect 14152 1180 14224 1214
rect 14452 1180 14524 1214
rect 14752 1180 14824 1214
rect 15052 1180 15124 1214
rect 15352 1180 15388 1214
rect 88 1168 15388 1180
rect 192 1130 284 1136
rect 192 1096 204 1130
rect 272 1096 284 1130
rect 192 1090 284 1096
rect 492 1130 584 1136
rect 492 1096 504 1130
rect 572 1096 584 1130
rect 492 1090 584 1096
rect 792 1130 884 1136
rect 792 1096 804 1130
rect 872 1096 884 1130
rect 792 1090 884 1096
rect 1092 1130 1184 1136
rect 1092 1096 1104 1130
rect 1172 1096 1184 1130
rect 1092 1090 1184 1096
rect 1392 1130 1484 1136
rect 1392 1096 1404 1130
rect 1472 1096 1484 1130
rect 1392 1090 1484 1096
rect 1692 1130 1784 1136
rect 1692 1096 1704 1130
rect 1772 1096 1784 1130
rect 1692 1090 1784 1096
rect 1992 1130 2084 1136
rect 1992 1096 2004 1130
rect 2072 1096 2084 1130
rect 1992 1090 2084 1096
rect 2292 1130 2384 1136
rect 2292 1096 2304 1130
rect 2372 1096 2384 1130
rect 2292 1090 2384 1096
rect 2592 1130 2684 1136
rect 2592 1096 2604 1130
rect 2672 1096 2684 1130
rect 2592 1090 2684 1096
rect 2892 1130 2984 1136
rect 2892 1096 2904 1130
rect 2972 1096 2984 1130
rect 2892 1090 2984 1096
rect 3192 1130 3284 1136
rect 3192 1096 3204 1130
rect 3272 1096 3284 1130
rect 3192 1090 3284 1096
rect 3492 1130 3584 1136
rect 3492 1096 3504 1130
rect 3572 1096 3584 1130
rect 3492 1090 3584 1096
rect 3792 1130 3884 1136
rect 3792 1096 3804 1130
rect 3872 1096 3884 1130
rect 3792 1090 3884 1096
rect 4092 1130 4184 1136
rect 4092 1096 4104 1130
rect 4172 1096 4184 1130
rect 4092 1090 4184 1096
rect 4392 1130 4484 1136
rect 4392 1096 4404 1130
rect 4472 1096 4484 1130
rect 4392 1090 4484 1096
rect 4692 1130 4784 1136
rect 4692 1096 4704 1130
rect 4772 1096 4784 1130
rect 4692 1090 4784 1096
rect 4992 1130 5084 1136
rect 4992 1096 5004 1130
rect 5072 1096 5084 1130
rect 4992 1090 5084 1096
rect 5292 1130 5384 1136
rect 5292 1096 5304 1130
rect 5372 1096 5384 1130
rect 5292 1090 5384 1096
rect 5592 1130 5684 1136
rect 5592 1096 5604 1130
rect 5672 1096 5684 1130
rect 5592 1090 5684 1096
rect 5892 1130 5984 1136
rect 5892 1096 5904 1130
rect 5972 1096 5984 1130
rect 5892 1090 5984 1096
rect 6192 1130 6284 1136
rect 6192 1096 6204 1130
rect 6272 1096 6284 1130
rect 6192 1090 6284 1096
rect 6492 1130 6584 1136
rect 6492 1096 6504 1130
rect 6572 1096 6584 1130
rect 6492 1090 6584 1096
rect 6792 1130 6884 1136
rect 6792 1096 6804 1130
rect 6872 1096 6884 1130
rect 6792 1090 6884 1096
rect 7092 1130 7184 1136
rect 7092 1096 7104 1130
rect 7172 1096 7184 1130
rect 7092 1090 7184 1096
rect 7392 1130 7484 1136
rect 7392 1096 7404 1130
rect 7472 1096 7484 1130
rect 7392 1090 7484 1096
rect 7692 1130 7784 1136
rect 7692 1096 7704 1130
rect 7772 1096 7784 1130
rect 7692 1090 7784 1096
rect 7992 1130 8084 1136
rect 7992 1096 8004 1130
rect 8072 1096 8084 1130
rect 7992 1090 8084 1096
rect 8292 1130 8384 1136
rect 8292 1096 8304 1130
rect 8372 1096 8384 1130
rect 8292 1090 8384 1096
rect 8592 1130 8684 1136
rect 8592 1096 8604 1130
rect 8672 1096 8684 1130
rect 8592 1090 8684 1096
rect 8892 1130 8984 1136
rect 8892 1096 8904 1130
rect 8972 1096 8984 1130
rect 8892 1090 8984 1096
rect 9192 1130 9284 1136
rect 9192 1096 9204 1130
rect 9272 1096 9284 1130
rect 9192 1090 9284 1096
rect 9492 1130 9584 1136
rect 9492 1096 9504 1130
rect 9572 1096 9584 1130
rect 9492 1090 9584 1096
rect 9792 1130 9884 1136
rect 9792 1096 9804 1130
rect 9872 1096 9884 1130
rect 9792 1090 9884 1096
rect 10092 1130 10184 1136
rect 10092 1096 10104 1130
rect 10172 1096 10184 1130
rect 10092 1090 10184 1096
rect 10392 1130 10484 1136
rect 10392 1096 10404 1130
rect 10472 1096 10484 1130
rect 10392 1090 10484 1096
rect 10692 1130 10784 1136
rect 10692 1096 10704 1130
rect 10772 1096 10784 1130
rect 10692 1090 10784 1096
rect 10992 1130 11084 1136
rect 10992 1096 11004 1130
rect 11072 1096 11084 1130
rect 10992 1090 11084 1096
rect 11292 1130 11384 1136
rect 11292 1096 11304 1130
rect 11372 1096 11384 1130
rect 11292 1090 11384 1096
rect 11592 1130 11684 1136
rect 11592 1096 11604 1130
rect 11672 1096 11684 1130
rect 11592 1090 11684 1096
rect 11892 1130 11984 1136
rect 11892 1096 11904 1130
rect 11972 1096 11984 1130
rect 11892 1090 11984 1096
rect 12192 1130 12284 1136
rect 12192 1096 12204 1130
rect 12272 1096 12284 1130
rect 12192 1090 12284 1096
rect 12492 1130 12584 1136
rect 12492 1096 12504 1130
rect 12572 1096 12584 1130
rect 12492 1090 12584 1096
rect 12792 1130 12884 1136
rect 12792 1096 12804 1130
rect 12872 1096 12884 1130
rect 12792 1090 12884 1096
rect 13092 1130 13184 1136
rect 13092 1096 13104 1130
rect 13172 1096 13184 1130
rect 13092 1090 13184 1096
rect 13392 1130 13484 1136
rect 13392 1096 13404 1130
rect 13472 1096 13484 1130
rect 13392 1090 13484 1096
rect 13692 1130 13784 1136
rect 13692 1096 13704 1130
rect 13772 1096 13784 1130
rect 13692 1090 13784 1096
rect 13992 1130 14084 1136
rect 13992 1096 14004 1130
rect 14072 1096 14084 1130
rect 13992 1090 14084 1096
rect 14292 1130 14384 1136
rect 14292 1096 14304 1130
rect 14372 1096 14384 1130
rect 14292 1090 14384 1096
rect 14592 1130 14684 1136
rect 14592 1096 14604 1130
rect 14672 1096 14684 1130
rect 14592 1090 14684 1096
rect 14892 1130 14984 1136
rect 14892 1096 14904 1130
rect 14972 1096 14984 1130
rect 14892 1090 14984 1096
rect 15192 1130 15284 1136
rect 15192 1096 15204 1130
rect 15272 1096 15284 1130
rect 15192 1090 15284 1096
rect 130 1049 164 1053
rect 124 1037 170 1049
rect 124 861 130 1037
rect 164 861 170 1037
rect 124 849 170 861
rect 130 845 164 849
rect 221 808 255 1090
rect 312 1049 346 1053
rect 430 1049 464 1053
rect 306 1037 352 1049
rect 306 861 312 1037
rect 346 861 352 1037
rect 306 849 352 861
rect 424 1037 470 1049
rect 424 861 430 1037
rect 464 861 470 1037
rect 424 849 470 861
rect 312 845 346 849
rect 430 845 464 849
rect 521 808 555 1090
rect 612 1049 646 1053
rect 730 1049 764 1053
rect 606 1037 652 1049
rect 606 861 612 1037
rect 646 861 652 1037
rect 606 849 652 861
rect 724 1037 770 1049
rect 724 861 730 1037
rect 764 861 770 1037
rect 724 849 770 861
rect 612 845 646 849
rect 730 845 764 849
rect 821 808 855 1090
rect 912 1049 946 1053
rect 1030 1049 1064 1053
rect 906 1037 952 1049
rect 906 861 912 1037
rect 946 861 952 1037
rect 906 849 952 861
rect 1024 1037 1070 1049
rect 1024 861 1030 1037
rect 1064 861 1070 1037
rect 1024 849 1070 861
rect 912 845 946 849
rect 1030 845 1064 849
rect 1121 808 1155 1090
rect 1212 1049 1246 1053
rect 1330 1049 1364 1053
rect 1206 1037 1252 1049
rect 1206 861 1212 1037
rect 1246 861 1252 1037
rect 1206 849 1252 861
rect 1324 1037 1370 1049
rect 1324 861 1330 1037
rect 1364 861 1370 1037
rect 1324 849 1370 861
rect 1212 845 1246 849
rect 1330 845 1364 849
rect 1421 808 1455 1090
rect 1512 1049 1546 1053
rect 1630 1049 1664 1053
rect 1506 1037 1552 1049
rect 1506 861 1512 1037
rect 1546 861 1552 1037
rect 1506 849 1552 861
rect 1624 1037 1670 1049
rect 1624 861 1630 1037
rect 1664 861 1670 1037
rect 1624 849 1670 861
rect 1512 845 1546 849
rect 1630 845 1664 849
rect 1721 808 1755 1090
rect 1812 1049 1846 1053
rect 1930 1049 1964 1053
rect 1806 1037 1852 1049
rect 1806 861 1812 1037
rect 1846 861 1852 1037
rect 1806 849 1852 861
rect 1924 1037 1970 1049
rect 1924 861 1930 1037
rect 1964 861 1970 1037
rect 1924 849 1970 861
rect 1812 845 1846 849
rect 1930 845 1964 849
rect 2021 808 2055 1090
rect 2112 1049 2146 1053
rect 2230 1049 2264 1053
rect 2106 1037 2152 1049
rect 2106 861 2112 1037
rect 2146 861 2152 1037
rect 2106 849 2152 861
rect 2224 1037 2270 1049
rect 2224 861 2230 1037
rect 2264 861 2270 1037
rect 2224 849 2270 861
rect 2112 845 2146 849
rect 2230 845 2264 849
rect 2321 808 2355 1090
rect 2412 1049 2446 1053
rect 2530 1049 2564 1053
rect 2406 1037 2452 1049
rect 2406 861 2412 1037
rect 2446 861 2452 1037
rect 2406 849 2452 861
rect 2524 1037 2570 1049
rect 2524 861 2530 1037
rect 2564 861 2570 1037
rect 2524 849 2570 861
rect 2412 845 2446 849
rect 2530 845 2564 849
rect 2621 808 2655 1090
rect 2712 1049 2746 1053
rect 2830 1049 2864 1053
rect 2706 1037 2752 1049
rect 2706 861 2712 1037
rect 2746 861 2752 1037
rect 2706 849 2752 861
rect 2824 1037 2870 1049
rect 2824 861 2830 1037
rect 2864 861 2870 1037
rect 2824 849 2870 861
rect 2712 845 2746 849
rect 2830 845 2864 849
rect 2921 808 2955 1090
rect 3012 1049 3046 1053
rect 3130 1049 3164 1053
rect 3006 1037 3052 1049
rect 3006 861 3012 1037
rect 3046 861 3052 1037
rect 3006 849 3052 861
rect 3124 1037 3170 1049
rect 3124 861 3130 1037
rect 3164 861 3170 1037
rect 3124 849 3170 861
rect 3012 845 3046 849
rect 3130 845 3164 849
rect 3221 808 3255 1090
rect 3312 1049 3346 1053
rect 3430 1049 3464 1053
rect 3306 1037 3352 1049
rect 3306 861 3312 1037
rect 3346 861 3352 1037
rect 3306 849 3352 861
rect 3424 1037 3470 1049
rect 3424 861 3430 1037
rect 3464 861 3470 1037
rect 3424 849 3470 861
rect 3312 845 3346 849
rect 3430 845 3464 849
rect 3521 808 3555 1090
rect 3612 1049 3646 1053
rect 3730 1049 3764 1053
rect 3606 1037 3652 1049
rect 3606 861 3612 1037
rect 3646 861 3652 1037
rect 3606 849 3652 861
rect 3724 1037 3770 1049
rect 3724 861 3730 1037
rect 3764 861 3770 1037
rect 3724 849 3770 861
rect 3612 845 3646 849
rect 3730 845 3764 849
rect 3821 808 3855 1090
rect 3912 1049 3946 1053
rect 4030 1049 4064 1053
rect 3906 1037 3952 1049
rect 3906 861 3912 1037
rect 3946 861 3952 1037
rect 3906 849 3952 861
rect 4024 1037 4070 1049
rect 4024 861 4030 1037
rect 4064 861 4070 1037
rect 4024 849 4070 861
rect 3912 845 3946 849
rect 4030 845 4064 849
rect 4121 808 4155 1090
rect 4212 1049 4246 1053
rect 4330 1049 4364 1053
rect 4206 1037 4252 1049
rect 4206 861 4212 1037
rect 4246 861 4252 1037
rect 4206 849 4252 861
rect 4324 1037 4370 1049
rect 4324 861 4330 1037
rect 4364 861 4370 1037
rect 4324 849 4370 861
rect 4212 845 4246 849
rect 4330 845 4364 849
rect 4421 808 4455 1090
rect 4512 1049 4546 1053
rect 4630 1049 4664 1053
rect 4506 1037 4552 1049
rect 4506 861 4512 1037
rect 4546 861 4552 1037
rect 4506 849 4552 861
rect 4624 1037 4670 1049
rect 4624 861 4630 1037
rect 4664 861 4670 1037
rect 4624 849 4670 861
rect 4512 845 4546 849
rect 4630 845 4664 849
rect 4721 808 4755 1090
rect 4812 1049 4846 1053
rect 4930 1049 4964 1053
rect 4806 1037 4852 1049
rect 4806 861 4812 1037
rect 4846 861 4852 1037
rect 4806 849 4852 861
rect 4924 1037 4970 1049
rect 4924 861 4930 1037
rect 4964 861 4970 1037
rect 4924 849 4970 861
rect 4812 845 4846 849
rect 4930 845 4964 849
rect 5021 808 5055 1090
rect 5112 1049 5146 1053
rect 5230 1049 5264 1053
rect 5106 1037 5152 1049
rect 5106 861 5112 1037
rect 5146 861 5152 1037
rect 5106 849 5152 861
rect 5224 1037 5270 1049
rect 5224 861 5230 1037
rect 5264 861 5270 1037
rect 5224 849 5270 861
rect 5112 845 5146 849
rect 5230 845 5264 849
rect 5321 808 5355 1090
rect 5412 1049 5446 1053
rect 5530 1049 5564 1053
rect 5406 1037 5452 1049
rect 5406 861 5412 1037
rect 5446 861 5452 1037
rect 5406 849 5452 861
rect 5524 1037 5570 1049
rect 5524 861 5530 1037
rect 5564 861 5570 1037
rect 5524 849 5570 861
rect 5412 845 5446 849
rect 5530 845 5564 849
rect 5621 808 5655 1090
rect 5712 1049 5746 1053
rect 5830 1049 5864 1053
rect 5706 1037 5752 1049
rect 5706 861 5712 1037
rect 5746 861 5752 1037
rect 5706 849 5752 861
rect 5824 1037 5870 1049
rect 5824 861 5830 1037
rect 5864 861 5870 1037
rect 5824 849 5870 861
rect 5712 845 5746 849
rect 5830 845 5864 849
rect 5921 808 5955 1090
rect 6012 1049 6046 1053
rect 6130 1049 6164 1053
rect 6006 1037 6052 1049
rect 6006 861 6012 1037
rect 6046 861 6052 1037
rect 6006 849 6052 861
rect 6124 1037 6170 1049
rect 6124 861 6130 1037
rect 6164 861 6170 1037
rect 6124 849 6170 861
rect 6012 845 6046 849
rect 6130 845 6164 849
rect 6221 808 6255 1090
rect 6312 1049 6346 1053
rect 6430 1049 6464 1053
rect 6306 1037 6352 1049
rect 6306 861 6312 1037
rect 6346 861 6352 1037
rect 6306 849 6352 861
rect 6424 1037 6470 1049
rect 6424 861 6430 1037
rect 6464 861 6470 1037
rect 6424 849 6470 861
rect 6312 845 6346 849
rect 6430 845 6464 849
rect 6521 808 6555 1090
rect 6612 1049 6646 1053
rect 6730 1049 6764 1053
rect 6606 1037 6652 1049
rect 6606 861 6612 1037
rect 6646 861 6652 1037
rect 6606 849 6652 861
rect 6724 1037 6770 1049
rect 6724 861 6730 1037
rect 6764 861 6770 1037
rect 6724 849 6770 861
rect 6612 845 6646 849
rect 6730 845 6764 849
rect 6821 808 6855 1090
rect 6912 1049 6946 1053
rect 7030 1049 7064 1053
rect 6906 1037 6952 1049
rect 6906 861 6912 1037
rect 6946 861 6952 1037
rect 6906 849 6952 861
rect 7024 1037 7070 1049
rect 7024 861 7030 1037
rect 7064 861 7070 1037
rect 7024 849 7070 861
rect 6912 845 6946 849
rect 7030 845 7064 849
rect 7121 808 7155 1090
rect 7212 1049 7246 1053
rect 7330 1049 7364 1053
rect 7206 1037 7252 1049
rect 7206 861 7212 1037
rect 7246 861 7252 1037
rect 7206 849 7252 861
rect 7324 1037 7370 1049
rect 7324 861 7330 1037
rect 7364 861 7370 1037
rect 7324 849 7370 861
rect 7212 845 7246 849
rect 7330 845 7364 849
rect 7421 808 7455 1090
rect 7512 1049 7546 1053
rect 7630 1049 7664 1053
rect 7506 1037 7552 1049
rect 7506 861 7512 1037
rect 7546 861 7552 1037
rect 7506 849 7552 861
rect 7624 1037 7670 1049
rect 7624 861 7630 1037
rect 7664 861 7670 1037
rect 7624 849 7670 861
rect 7512 845 7546 849
rect 7630 845 7664 849
rect 7721 808 7755 1090
rect 7812 1049 7846 1053
rect 7930 1049 7964 1053
rect 7806 1037 7852 1049
rect 7806 861 7812 1037
rect 7846 861 7852 1037
rect 7806 849 7852 861
rect 7924 1037 7970 1049
rect 7924 861 7930 1037
rect 7964 861 7970 1037
rect 7924 849 7970 861
rect 7812 845 7846 849
rect 7930 845 7964 849
rect 8021 808 8055 1090
rect 8112 1049 8146 1053
rect 8230 1049 8264 1053
rect 8106 1037 8152 1049
rect 8106 861 8112 1037
rect 8146 861 8152 1037
rect 8106 849 8152 861
rect 8224 1037 8270 1049
rect 8224 861 8230 1037
rect 8264 861 8270 1037
rect 8224 849 8270 861
rect 8112 845 8146 849
rect 8230 845 8264 849
rect 8321 808 8355 1090
rect 8412 1049 8446 1053
rect 8530 1049 8564 1053
rect 8406 1037 8452 1049
rect 8406 861 8412 1037
rect 8446 861 8452 1037
rect 8406 849 8452 861
rect 8524 1037 8570 1049
rect 8524 861 8530 1037
rect 8564 861 8570 1037
rect 8524 849 8570 861
rect 8412 845 8446 849
rect 8530 845 8564 849
rect 8621 808 8655 1090
rect 8712 1049 8746 1053
rect 8830 1049 8864 1053
rect 8706 1037 8752 1049
rect 8706 861 8712 1037
rect 8746 861 8752 1037
rect 8706 849 8752 861
rect 8824 1037 8870 1049
rect 8824 861 8830 1037
rect 8864 861 8870 1037
rect 8824 849 8870 861
rect 8712 845 8746 849
rect 8830 845 8864 849
rect 8921 808 8955 1090
rect 9012 1049 9046 1053
rect 9130 1049 9164 1053
rect 9006 1037 9052 1049
rect 9006 861 9012 1037
rect 9046 861 9052 1037
rect 9006 849 9052 861
rect 9124 1037 9170 1049
rect 9124 861 9130 1037
rect 9164 861 9170 1037
rect 9124 849 9170 861
rect 9012 845 9046 849
rect 9130 845 9164 849
rect 9221 808 9255 1090
rect 9312 1049 9346 1053
rect 9430 1049 9464 1053
rect 9306 1037 9352 1049
rect 9306 861 9312 1037
rect 9346 861 9352 1037
rect 9306 849 9352 861
rect 9424 1037 9470 1049
rect 9424 861 9430 1037
rect 9464 861 9470 1037
rect 9424 849 9470 861
rect 9312 845 9346 849
rect 9430 845 9464 849
rect 9521 808 9555 1090
rect 9612 1049 9646 1053
rect 9730 1049 9764 1053
rect 9606 1037 9652 1049
rect 9606 861 9612 1037
rect 9646 861 9652 1037
rect 9606 849 9652 861
rect 9724 1037 9770 1049
rect 9724 861 9730 1037
rect 9764 861 9770 1037
rect 9724 849 9770 861
rect 9612 845 9646 849
rect 9730 845 9764 849
rect 9821 808 9855 1090
rect 9912 1049 9946 1053
rect 10030 1049 10064 1053
rect 9906 1037 9952 1049
rect 9906 861 9912 1037
rect 9946 861 9952 1037
rect 9906 849 9952 861
rect 10024 1037 10070 1049
rect 10024 861 10030 1037
rect 10064 861 10070 1037
rect 10024 849 10070 861
rect 9912 845 9946 849
rect 10030 845 10064 849
rect 10121 808 10155 1090
rect 10212 1049 10246 1053
rect 10330 1049 10364 1053
rect 10206 1037 10252 1049
rect 10206 861 10212 1037
rect 10246 861 10252 1037
rect 10206 849 10252 861
rect 10324 1037 10370 1049
rect 10324 861 10330 1037
rect 10364 861 10370 1037
rect 10324 849 10370 861
rect 10212 845 10246 849
rect 10330 845 10364 849
rect 10421 808 10455 1090
rect 10512 1049 10546 1053
rect 10630 1049 10664 1053
rect 10506 1037 10552 1049
rect 10506 861 10512 1037
rect 10546 861 10552 1037
rect 10506 849 10552 861
rect 10624 1037 10670 1049
rect 10624 861 10630 1037
rect 10664 861 10670 1037
rect 10624 849 10670 861
rect 10512 845 10546 849
rect 10630 845 10664 849
rect 10721 808 10755 1090
rect 10812 1049 10846 1053
rect 10930 1049 10964 1053
rect 10806 1037 10852 1049
rect 10806 861 10812 1037
rect 10846 861 10852 1037
rect 10806 849 10852 861
rect 10924 1037 10970 1049
rect 10924 861 10930 1037
rect 10964 861 10970 1037
rect 10924 849 10970 861
rect 10812 845 10846 849
rect 10930 845 10964 849
rect 11021 808 11055 1090
rect 11112 1049 11146 1053
rect 11230 1049 11264 1053
rect 11106 1037 11152 1049
rect 11106 861 11112 1037
rect 11146 861 11152 1037
rect 11106 849 11152 861
rect 11224 1037 11270 1049
rect 11224 861 11230 1037
rect 11264 861 11270 1037
rect 11224 849 11270 861
rect 11112 845 11146 849
rect 11230 845 11264 849
rect 11321 808 11355 1090
rect 11412 1049 11446 1053
rect 11530 1049 11564 1053
rect 11406 1037 11452 1049
rect 11406 861 11412 1037
rect 11446 861 11452 1037
rect 11406 849 11452 861
rect 11524 1037 11570 1049
rect 11524 861 11530 1037
rect 11564 861 11570 1037
rect 11524 849 11570 861
rect 11412 845 11446 849
rect 11530 845 11564 849
rect 11621 808 11655 1090
rect 11712 1049 11746 1053
rect 11830 1049 11864 1053
rect 11706 1037 11752 1049
rect 11706 861 11712 1037
rect 11746 861 11752 1037
rect 11706 849 11752 861
rect 11824 1037 11870 1049
rect 11824 861 11830 1037
rect 11864 861 11870 1037
rect 11824 849 11870 861
rect 11712 845 11746 849
rect 11830 845 11864 849
rect 11921 808 11955 1090
rect 12012 1049 12046 1053
rect 12130 1049 12164 1053
rect 12006 1037 12052 1049
rect 12006 861 12012 1037
rect 12046 861 12052 1037
rect 12006 849 12052 861
rect 12124 1037 12170 1049
rect 12124 861 12130 1037
rect 12164 861 12170 1037
rect 12124 849 12170 861
rect 12012 845 12046 849
rect 12130 845 12164 849
rect 12221 808 12255 1090
rect 12312 1049 12346 1053
rect 12430 1049 12464 1053
rect 12306 1037 12352 1049
rect 12306 861 12312 1037
rect 12346 861 12352 1037
rect 12306 849 12352 861
rect 12424 1037 12470 1049
rect 12424 861 12430 1037
rect 12464 861 12470 1037
rect 12424 849 12470 861
rect 12312 845 12346 849
rect 12430 845 12464 849
rect 12521 808 12555 1090
rect 12612 1049 12646 1053
rect 12730 1049 12764 1053
rect 12606 1037 12652 1049
rect 12606 861 12612 1037
rect 12646 861 12652 1037
rect 12606 849 12652 861
rect 12724 1037 12770 1049
rect 12724 861 12730 1037
rect 12764 861 12770 1037
rect 12724 849 12770 861
rect 12612 845 12646 849
rect 12730 845 12764 849
rect 12821 808 12855 1090
rect 12912 1049 12946 1053
rect 13030 1049 13064 1053
rect 12906 1037 12952 1049
rect 12906 861 12912 1037
rect 12946 861 12952 1037
rect 12906 849 12952 861
rect 13024 1037 13070 1049
rect 13024 861 13030 1037
rect 13064 861 13070 1037
rect 13024 849 13070 861
rect 12912 845 12946 849
rect 13030 845 13064 849
rect 13121 808 13155 1090
rect 13212 1049 13246 1053
rect 13330 1049 13364 1053
rect 13206 1037 13252 1049
rect 13206 861 13212 1037
rect 13246 861 13252 1037
rect 13206 849 13252 861
rect 13324 1037 13370 1049
rect 13324 861 13330 1037
rect 13364 861 13370 1037
rect 13324 849 13370 861
rect 13212 845 13246 849
rect 13330 845 13364 849
rect 13421 808 13455 1090
rect 13512 1049 13546 1053
rect 13630 1049 13664 1053
rect 13506 1037 13552 1049
rect 13506 861 13512 1037
rect 13546 861 13552 1037
rect 13506 849 13552 861
rect 13624 1037 13670 1049
rect 13624 861 13630 1037
rect 13664 861 13670 1037
rect 13624 849 13670 861
rect 13512 845 13546 849
rect 13630 845 13664 849
rect 13721 808 13755 1090
rect 13812 1049 13846 1053
rect 13930 1049 13964 1053
rect 13806 1037 13852 1049
rect 13806 861 13812 1037
rect 13846 861 13852 1037
rect 13806 849 13852 861
rect 13924 1037 13970 1049
rect 13924 861 13930 1037
rect 13964 861 13970 1037
rect 13924 849 13970 861
rect 13812 845 13846 849
rect 13930 845 13964 849
rect 14021 808 14055 1090
rect 14112 1049 14146 1053
rect 14230 1049 14264 1053
rect 14106 1037 14152 1049
rect 14106 861 14112 1037
rect 14146 861 14152 1037
rect 14106 849 14152 861
rect 14224 1037 14270 1049
rect 14224 861 14230 1037
rect 14264 861 14270 1037
rect 14224 849 14270 861
rect 14112 845 14146 849
rect 14230 845 14264 849
rect 14321 808 14355 1090
rect 14412 1049 14446 1053
rect 14530 1049 14564 1053
rect 14406 1037 14452 1049
rect 14406 861 14412 1037
rect 14446 861 14452 1037
rect 14406 849 14452 861
rect 14524 1037 14570 1049
rect 14524 861 14530 1037
rect 14564 861 14570 1037
rect 14524 849 14570 861
rect 14412 845 14446 849
rect 14530 845 14564 849
rect 14621 808 14655 1090
rect 14712 1049 14746 1053
rect 14830 1049 14864 1053
rect 14706 1037 14752 1049
rect 14706 861 14712 1037
rect 14746 861 14752 1037
rect 14706 849 14752 861
rect 14824 1037 14870 1049
rect 14824 861 14830 1037
rect 14864 861 14870 1037
rect 14824 849 14870 861
rect 14712 845 14746 849
rect 14830 845 14864 849
rect 14921 808 14955 1090
rect 15012 1049 15046 1053
rect 15130 1049 15164 1053
rect 15006 1037 15052 1049
rect 15006 861 15012 1037
rect 15046 861 15052 1037
rect 15006 849 15052 861
rect 15124 1037 15170 1049
rect 15124 861 15130 1037
rect 15164 861 15170 1037
rect 15124 849 15170 861
rect 15012 845 15046 849
rect 15130 845 15164 849
rect 15221 808 15255 1090
rect 15312 1049 15346 1053
rect 15306 1037 15352 1049
rect 15306 861 15312 1037
rect 15346 861 15352 1037
rect 15306 849 15352 861
rect 15312 845 15346 849
rect 192 802 284 808
rect 192 768 204 802
rect 272 768 284 802
rect 192 762 284 768
rect 492 802 584 808
rect 492 768 504 802
rect 572 768 584 802
rect 492 762 584 768
rect 792 802 884 808
rect 792 768 804 802
rect 872 768 884 802
rect 792 762 884 768
rect 1092 802 1184 808
rect 1092 768 1104 802
rect 1172 768 1184 802
rect 1092 762 1184 768
rect 1392 802 1484 808
rect 1392 768 1404 802
rect 1472 768 1484 802
rect 1392 762 1484 768
rect 1692 802 1784 808
rect 1692 768 1704 802
rect 1772 768 1784 802
rect 1692 762 1784 768
rect 1992 802 2084 808
rect 1992 768 2004 802
rect 2072 768 2084 802
rect 1992 762 2084 768
rect 2292 802 2384 808
rect 2292 768 2304 802
rect 2372 768 2384 802
rect 2292 762 2384 768
rect 2592 802 2684 808
rect 2592 768 2604 802
rect 2672 768 2684 802
rect 2592 762 2684 768
rect 2892 802 2984 808
rect 2892 768 2904 802
rect 2972 768 2984 802
rect 2892 762 2984 768
rect 3192 802 3284 808
rect 3192 768 3204 802
rect 3272 768 3284 802
rect 3192 762 3284 768
rect 3492 802 3584 808
rect 3492 768 3504 802
rect 3572 768 3584 802
rect 3492 762 3584 768
rect 3792 802 3884 808
rect 3792 768 3804 802
rect 3872 768 3884 802
rect 3792 762 3884 768
rect 4092 802 4184 808
rect 4092 768 4104 802
rect 4172 768 4184 802
rect 4092 762 4184 768
rect 4392 802 4484 808
rect 4392 768 4404 802
rect 4472 768 4484 802
rect 4392 762 4484 768
rect 4692 802 4784 808
rect 4692 768 4704 802
rect 4772 768 4784 802
rect 4692 762 4784 768
rect 4992 802 5084 808
rect 4992 768 5004 802
rect 5072 768 5084 802
rect 4992 762 5084 768
rect 5292 802 5384 808
rect 5292 768 5304 802
rect 5372 768 5384 802
rect 5292 762 5384 768
rect 5592 802 5684 808
rect 5592 768 5604 802
rect 5672 768 5684 802
rect 5592 762 5684 768
rect 5892 802 5984 808
rect 5892 768 5904 802
rect 5972 768 5984 802
rect 5892 762 5984 768
rect 6192 802 6284 808
rect 6192 768 6204 802
rect 6272 768 6284 802
rect 6192 762 6284 768
rect 6492 802 6584 808
rect 6492 768 6504 802
rect 6572 768 6584 802
rect 6492 762 6584 768
rect 6792 802 6884 808
rect 6792 768 6804 802
rect 6872 768 6884 802
rect 6792 762 6884 768
rect 7092 802 7184 808
rect 7092 768 7104 802
rect 7172 768 7184 802
rect 7092 762 7184 768
rect 7392 802 7484 808
rect 7392 768 7404 802
rect 7472 768 7484 802
rect 7392 762 7484 768
rect 7692 802 7784 808
rect 7692 768 7704 802
rect 7772 768 7784 802
rect 7692 762 7784 768
rect 7992 802 8084 808
rect 7992 768 8004 802
rect 8072 768 8084 802
rect 7992 762 8084 768
rect 8292 802 8384 808
rect 8292 768 8304 802
rect 8372 768 8384 802
rect 8292 762 8384 768
rect 8592 802 8684 808
rect 8592 768 8604 802
rect 8672 768 8684 802
rect 8592 762 8684 768
rect 8892 802 8984 808
rect 8892 768 8904 802
rect 8972 768 8984 802
rect 8892 762 8984 768
rect 9192 802 9284 808
rect 9192 768 9204 802
rect 9272 768 9284 802
rect 9192 762 9284 768
rect 9492 802 9584 808
rect 9492 768 9504 802
rect 9572 768 9584 802
rect 9492 762 9584 768
rect 9792 802 9884 808
rect 9792 768 9804 802
rect 9872 768 9884 802
rect 9792 762 9884 768
rect 10092 802 10184 808
rect 10092 768 10104 802
rect 10172 768 10184 802
rect 10092 762 10184 768
rect 10392 802 10484 808
rect 10392 768 10404 802
rect 10472 768 10484 802
rect 10392 762 10484 768
rect 10692 802 10784 808
rect 10692 768 10704 802
rect 10772 768 10784 802
rect 10692 762 10784 768
rect 10992 802 11084 808
rect 10992 768 11004 802
rect 11072 768 11084 802
rect 10992 762 11084 768
rect 11292 802 11384 808
rect 11292 768 11304 802
rect 11372 768 11384 802
rect 11292 762 11384 768
rect 11592 802 11684 808
rect 11592 768 11604 802
rect 11672 768 11684 802
rect 11592 762 11684 768
rect 11892 802 11984 808
rect 11892 768 11904 802
rect 11972 768 11984 802
rect 11892 762 11984 768
rect 12192 802 12284 808
rect 12192 768 12204 802
rect 12272 768 12284 802
rect 12192 762 12284 768
rect 12492 802 12584 808
rect 12492 768 12504 802
rect 12572 768 12584 802
rect 12492 762 12584 768
rect 12792 802 12884 808
rect 12792 768 12804 802
rect 12872 768 12884 802
rect 12792 762 12884 768
rect 13092 802 13184 808
rect 13092 768 13104 802
rect 13172 768 13184 802
rect 13092 762 13184 768
rect 13392 802 13484 808
rect 13392 768 13404 802
rect 13472 768 13484 802
rect 13392 762 13484 768
rect 13692 802 13784 808
rect 13692 768 13704 802
rect 13772 768 13784 802
rect 13692 762 13784 768
rect 13992 802 14084 808
rect 13992 768 14004 802
rect 14072 768 14084 802
rect 13992 762 14084 768
rect 14292 802 14384 808
rect 14292 768 14304 802
rect 14372 768 14384 802
rect 14292 762 14384 768
rect 14592 802 14684 808
rect 14592 768 14604 802
rect 14672 768 14684 802
rect 14592 762 14684 768
rect 14892 802 14984 808
rect 14892 768 14904 802
rect 14972 768 14984 802
rect 14892 762 14984 768
rect 15192 802 15284 808
rect 15192 768 15204 802
rect 15272 768 15284 802
rect 15192 762 15284 768
rect 192 415 284 421
rect 192 381 204 415
rect 272 381 284 415
rect 192 375 284 381
rect 492 415 584 421
rect 492 381 504 415
rect 572 381 584 415
rect 492 375 584 381
rect 792 415 884 421
rect 792 381 804 415
rect 872 381 884 415
rect 792 375 884 381
rect 1092 415 1184 421
rect 1092 381 1104 415
rect 1172 381 1184 415
rect 1092 375 1184 381
rect 1392 415 1484 421
rect 1392 381 1404 415
rect 1472 381 1484 415
rect 1392 375 1484 381
rect 1692 415 1784 421
rect 1692 381 1704 415
rect 1772 381 1784 415
rect 1692 375 1784 381
rect 1992 415 2084 421
rect 1992 381 2004 415
rect 2072 381 2084 415
rect 1992 375 2084 381
rect 2292 415 2384 421
rect 2292 381 2304 415
rect 2372 381 2384 415
rect 2292 375 2384 381
rect 2592 415 2684 421
rect 2592 381 2604 415
rect 2672 381 2684 415
rect 2592 375 2684 381
rect 2892 415 2984 421
rect 2892 381 2904 415
rect 2972 381 2984 415
rect 2892 375 2984 381
rect 3192 415 3284 421
rect 3192 381 3204 415
rect 3272 381 3284 415
rect 3192 375 3284 381
rect 3492 415 3584 421
rect 3492 381 3504 415
rect 3572 381 3584 415
rect 3492 375 3584 381
rect 3792 415 3884 421
rect 3792 381 3804 415
rect 3872 381 3884 415
rect 3792 375 3884 381
rect 4092 415 4184 421
rect 4092 381 4104 415
rect 4172 381 4184 415
rect 4092 375 4184 381
rect 4392 415 4484 421
rect 4392 381 4404 415
rect 4472 381 4484 415
rect 4392 375 4484 381
rect 4692 415 4784 421
rect 4692 381 4704 415
rect 4772 381 4784 415
rect 4692 375 4784 381
rect 4992 415 5084 421
rect 4992 381 5004 415
rect 5072 381 5084 415
rect 4992 375 5084 381
rect 5292 415 5384 421
rect 5292 381 5304 415
rect 5372 381 5384 415
rect 5292 375 5384 381
rect 5592 415 5684 421
rect 5592 381 5604 415
rect 5672 381 5684 415
rect 5592 375 5684 381
rect 5892 415 5984 421
rect 5892 381 5904 415
rect 5972 381 5984 415
rect 5892 375 5984 381
rect 6192 415 6284 421
rect 6192 381 6204 415
rect 6272 381 6284 415
rect 6192 375 6284 381
rect 6492 415 6584 421
rect 6492 381 6504 415
rect 6572 381 6584 415
rect 6492 375 6584 381
rect 6792 415 6884 421
rect 6792 381 6804 415
rect 6872 381 6884 415
rect 6792 375 6884 381
rect 7092 415 7184 421
rect 7092 381 7104 415
rect 7172 381 7184 415
rect 7092 375 7184 381
rect 7392 415 7484 421
rect 7392 381 7404 415
rect 7472 381 7484 415
rect 7392 375 7484 381
rect 7692 415 7784 421
rect 7692 381 7704 415
rect 7772 381 7784 415
rect 7692 375 7784 381
rect 7992 415 8084 421
rect 7992 381 8004 415
rect 8072 381 8084 415
rect 7992 375 8084 381
rect 8292 415 8384 421
rect 8292 381 8304 415
rect 8372 381 8384 415
rect 8292 375 8384 381
rect 8592 415 8684 421
rect 8592 381 8604 415
rect 8672 381 8684 415
rect 8592 375 8684 381
rect 8892 415 8984 421
rect 8892 381 8904 415
rect 8972 381 8984 415
rect 8892 375 8984 381
rect 9192 415 9284 421
rect 9192 381 9204 415
rect 9272 381 9284 415
rect 9192 375 9284 381
rect 9492 415 9584 421
rect 9492 381 9504 415
rect 9572 381 9584 415
rect 9492 375 9584 381
rect 9792 415 9884 421
rect 9792 381 9804 415
rect 9872 381 9884 415
rect 9792 375 9884 381
rect 10092 415 10184 421
rect 10092 381 10104 415
rect 10172 381 10184 415
rect 10092 375 10184 381
rect 10392 415 10484 421
rect 10392 381 10404 415
rect 10472 381 10484 415
rect 10392 375 10484 381
rect 10692 415 10784 421
rect 10692 381 10704 415
rect 10772 381 10784 415
rect 10692 375 10784 381
rect 10992 415 11084 421
rect 10992 381 11004 415
rect 11072 381 11084 415
rect 10992 375 11084 381
rect 11292 415 11384 421
rect 11292 381 11304 415
rect 11372 381 11384 415
rect 11292 375 11384 381
rect 11592 415 11684 421
rect 11592 381 11604 415
rect 11672 381 11684 415
rect 11592 375 11684 381
rect 11892 415 11984 421
rect 11892 381 11904 415
rect 11972 381 11984 415
rect 11892 375 11984 381
rect 12192 415 12284 421
rect 12192 381 12204 415
rect 12272 381 12284 415
rect 12192 375 12284 381
rect 12492 415 12584 421
rect 12492 381 12504 415
rect 12572 381 12584 415
rect 12492 375 12584 381
rect 12792 415 12884 421
rect 12792 381 12804 415
rect 12872 381 12884 415
rect 12792 375 12884 381
rect 13092 415 13184 421
rect 13092 381 13104 415
rect 13172 381 13184 415
rect 13092 375 13184 381
rect 13392 415 13484 421
rect 13392 381 13404 415
rect 13472 381 13484 415
rect 13392 375 13484 381
rect 13692 415 13784 421
rect 13692 381 13704 415
rect 13772 381 13784 415
rect 13692 375 13784 381
rect 13992 415 14084 421
rect 13992 381 14004 415
rect 14072 381 14084 415
rect 13992 375 14084 381
rect 14292 415 14384 421
rect 14292 381 14304 415
rect 14372 381 14384 415
rect 14292 375 14384 381
rect 14592 415 14684 421
rect 14592 381 14604 415
rect 14672 381 14684 415
rect 14592 375 14684 381
rect 14892 415 14984 421
rect 14892 381 14904 415
rect 14972 381 14984 415
rect 14892 375 14984 381
rect 15192 415 15284 421
rect 15192 381 15204 415
rect 15272 381 15284 415
rect 15192 375 15284 381
rect 130 343 164 347
rect 124 331 170 343
rect 124 225 130 331
rect 164 225 170 331
rect 124 213 170 225
rect 130 209 164 213
rect 221 181 255 375
rect 312 343 346 347
rect 430 343 464 347
rect 306 331 352 343
rect 306 225 312 331
rect 346 225 352 331
rect 306 213 352 225
rect 424 331 470 343
rect 424 225 430 331
rect 464 225 470 331
rect 424 213 470 225
rect 312 209 346 213
rect 430 209 464 213
rect 521 181 555 375
rect 612 343 646 347
rect 730 343 764 347
rect 606 331 652 343
rect 606 225 612 331
rect 646 225 652 331
rect 606 213 652 225
rect 724 331 770 343
rect 724 225 730 331
rect 764 225 770 331
rect 724 213 770 225
rect 612 209 646 213
rect 730 209 764 213
rect 821 181 855 375
rect 912 343 946 347
rect 1030 343 1064 347
rect 906 331 952 343
rect 906 225 912 331
rect 946 225 952 331
rect 906 213 952 225
rect 1024 331 1070 343
rect 1024 225 1030 331
rect 1064 225 1070 331
rect 1024 213 1070 225
rect 912 209 946 213
rect 1030 209 1064 213
rect 1121 181 1155 375
rect 1212 343 1246 347
rect 1330 343 1364 347
rect 1206 331 1252 343
rect 1206 225 1212 331
rect 1246 225 1252 331
rect 1206 213 1252 225
rect 1324 331 1370 343
rect 1324 225 1330 331
rect 1364 225 1370 331
rect 1324 213 1370 225
rect 1212 209 1246 213
rect 1330 209 1364 213
rect 1421 181 1455 375
rect 1512 343 1546 347
rect 1630 343 1664 347
rect 1506 331 1552 343
rect 1506 225 1512 331
rect 1546 225 1552 331
rect 1506 213 1552 225
rect 1624 331 1670 343
rect 1624 225 1630 331
rect 1664 225 1670 331
rect 1624 213 1670 225
rect 1512 209 1546 213
rect 1630 209 1664 213
rect 1721 181 1755 375
rect 1812 343 1846 347
rect 1930 343 1964 347
rect 1806 331 1852 343
rect 1806 225 1812 331
rect 1846 225 1852 331
rect 1806 213 1852 225
rect 1924 331 1970 343
rect 1924 225 1930 331
rect 1964 225 1970 331
rect 1924 213 1970 225
rect 1812 209 1846 213
rect 1930 209 1964 213
rect 2021 181 2055 375
rect 2112 343 2146 347
rect 2230 343 2264 347
rect 2106 331 2152 343
rect 2106 225 2112 331
rect 2146 225 2152 331
rect 2106 213 2152 225
rect 2224 331 2270 343
rect 2224 225 2230 331
rect 2264 225 2270 331
rect 2224 213 2270 225
rect 2112 209 2146 213
rect 2230 209 2264 213
rect 2321 181 2355 375
rect 2412 343 2446 347
rect 2530 343 2564 347
rect 2406 331 2452 343
rect 2406 225 2412 331
rect 2446 225 2452 331
rect 2406 213 2452 225
rect 2524 331 2570 343
rect 2524 225 2530 331
rect 2564 225 2570 331
rect 2524 213 2570 225
rect 2412 209 2446 213
rect 2530 209 2564 213
rect 2621 181 2655 375
rect 2712 343 2746 347
rect 2830 343 2864 347
rect 2706 331 2752 343
rect 2706 225 2712 331
rect 2746 225 2752 331
rect 2706 213 2752 225
rect 2824 331 2870 343
rect 2824 225 2830 331
rect 2864 225 2870 331
rect 2824 213 2870 225
rect 2712 209 2746 213
rect 2830 209 2864 213
rect 2921 181 2955 375
rect 3012 343 3046 347
rect 3130 343 3164 347
rect 3006 331 3052 343
rect 3006 225 3012 331
rect 3046 225 3052 331
rect 3006 213 3052 225
rect 3124 331 3170 343
rect 3124 225 3130 331
rect 3164 225 3170 331
rect 3124 213 3170 225
rect 3012 209 3046 213
rect 3130 209 3164 213
rect 3221 181 3255 375
rect 3312 343 3346 347
rect 3430 343 3464 347
rect 3306 331 3352 343
rect 3306 225 3312 331
rect 3346 225 3352 331
rect 3306 213 3352 225
rect 3424 331 3470 343
rect 3424 225 3430 331
rect 3464 225 3470 331
rect 3424 213 3470 225
rect 3312 209 3346 213
rect 3430 209 3464 213
rect 3521 181 3555 375
rect 3612 343 3646 347
rect 3730 343 3764 347
rect 3606 331 3652 343
rect 3606 225 3612 331
rect 3646 225 3652 331
rect 3606 213 3652 225
rect 3724 331 3770 343
rect 3724 225 3730 331
rect 3764 225 3770 331
rect 3724 213 3770 225
rect 3612 209 3646 213
rect 3730 209 3764 213
rect 3821 181 3855 375
rect 3912 343 3946 347
rect 4030 343 4064 347
rect 3906 331 3952 343
rect 3906 225 3912 331
rect 3946 225 3952 331
rect 3906 213 3952 225
rect 4024 331 4070 343
rect 4024 225 4030 331
rect 4064 225 4070 331
rect 4024 213 4070 225
rect 3912 209 3946 213
rect 4030 209 4064 213
rect 4121 181 4155 375
rect 4212 343 4246 347
rect 4330 343 4364 347
rect 4206 331 4252 343
rect 4206 225 4212 331
rect 4246 225 4252 331
rect 4206 213 4252 225
rect 4324 331 4370 343
rect 4324 225 4330 331
rect 4364 225 4370 331
rect 4324 213 4370 225
rect 4212 209 4246 213
rect 4330 209 4364 213
rect 4421 181 4455 375
rect 4512 343 4546 347
rect 4630 343 4664 347
rect 4506 331 4552 343
rect 4506 225 4512 331
rect 4546 225 4552 331
rect 4506 213 4552 225
rect 4624 331 4670 343
rect 4624 225 4630 331
rect 4664 225 4670 331
rect 4624 213 4670 225
rect 4512 209 4546 213
rect 4630 209 4664 213
rect 4721 181 4755 375
rect 4812 343 4846 347
rect 4930 343 4964 347
rect 4806 331 4852 343
rect 4806 225 4812 331
rect 4846 225 4852 331
rect 4806 213 4852 225
rect 4924 331 4970 343
rect 4924 225 4930 331
rect 4964 225 4970 331
rect 4924 213 4970 225
rect 4812 209 4846 213
rect 4930 209 4964 213
rect 5021 181 5055 375
rect 5112 343 5146 347
rect 5230 343 5264 347
rect 5106 331 5152 343
rect 5106 225 5112 331
rect 5146 225 5152 331
rect 5106 213 5152 225
rect 5224 331 5270 343
rect 5224 225 5230 331
rect 5264 225 5270 331
rect 5224 213 5270 225
rect 5112 209 5146 213
rect 5230 209 5264 213
rect 5321 181 5355 375
rect 5412 343 5446 347
rect 5530 343 5564 347
rect 5406 331 5452 343
rect 5406 225 5412 331
rect 5446 225 5452 331
rect 5406 213 5452 225
rect 5524 331 5570 343
rect 5524 225 5530 331
rect 5564 225 5570 331
rect 5524 213 5570 225
rect 5412 209 5446 213
rect 5530 209 5564 213
rect 5621 181 5655 375
rect 5712 343 5746 347
rect 5830 343 5864 347
rect 5706 331 5752 343
rect 5706 225 5712 331
rect 5746 225 5752 331
rect 5706 213 5752 225
rect 5824 331 5870 343
rect 5824 225 5830 331
rect 5864 225 5870 331
rect 5824 213 5870 225
rect 5712 209 5746 213
rect 5830 209 5864 213
rect 5921 181 5955 375
rect 6012 343 6046 347
rect 6130 343 6164 347
rect 6006 331 6052 343
rect 6006 225 6012 331
rect 6046 225 6052 331
rect 6006 213 6052 225
rect 6124 331 6170 343
rect 6124 225 6130 331
rect 6164 225 6170 331
rect 6124 213 6170 225
rect 6012 209 6046 213
rect 6130 209 6164 213
rect 6221 181 6255 375
rect 6312 343 6346 347
rect 6430 343 6464 347
rect 6306 331 6352 343
rect 6306 225 6312 331
rect 6346 225 6352 331
rect 6306 213 6352 225
rect 6424 331 6470 343
rect 6424 225 6430 331
rect 6464 225 6470 331
rect 6424 213 6470 225
rect 6312 209 6346 213
rect 6430 209 6464 213
rect 6521 181 6555 375
rect 6612 343 6646 347
rect 6730 343 6764 347
rect 6606 331 6652 343
rect 6606 225 6612 331
rect 6646 225 6652 331
rect 6606 213 6652 225
rect 6724 331 6770 343
rect 6724 225 6730 331
rect 6764 225 6770 331
rect 6724 213 6770 225
rect 6612 209 6646 213
rect 6730 209 6764 213
rect 6821 181 6855 375
rect 6912 343 6946 347
rect 7030 343 7064 347
rect 6906 331 6952 343
rect 6906 225 6912 331
rect 6946 225 6952 331
rect 6906 213 6952 225
rect 7024 331 7070 343
rect 7024 225 7030 331
rect 7064 225 7070 331
rect 7024 213 7070 225
rect 6912 209 6946 213
rect 7030 209 7064 213
rect 7121 181 7155 375
rect 7212 343 7246 347
rect 7330 343 7364 347
rect 7206 331 7252 343
rect 7206 225 7212 331
rect 7246 225 7252 331
rect 7206 213 7252 225
rect 7324 331 7370 343
rect 7324 225 7330 331
rect 7364 225 7370 331
rect 7324 213 7370 225
rect 7212 209 7246 213
rect 7330 209 7364 213
rect 7421 181 7455 375
rect 7512 343 7546 347
rect 7630 343 7664 347
rect 7506 331 7552 343
rect 7506 225 7512 331
rect 7546 225 7552 331
rect 7506 213 7552 225
rect 7624 331 7670 343
rect 7624 225 7630 331
rect 7664 225 7670 331
rect 7624 213 7670 225
rect 7512 209 7546 213
rect 7630 209 7664 213
rect 7721 181 7755 375
rect 7812 343 7846 347
rect 7930 343 7964 347
rect 7806 331 7852 343
rect 7806 225 7812 331
rect 7846 225 7852 331
rect 7806 213 7852 225
rect 7924 331 7970 343
rect 7924 225 7930 331
rect 7964 225 7970 331
rect 7924 213 7970 225
rect 7812 209 7846 213
rect 7930 209 7964 213
rect 8021 181 8055 375
rect 8112 343 8146 347
rect 8230 343 8264 347
rect 8106 331 8152 343
rect 8106 225 8112 331
rect 8146 225 8152 331
rect 8106 213 8152 225
rect 8224 331 8270 343
rect 8224 225 8230 331
rect 8264 225 8270 331
rect 8224 213 8270 225
rect 8112 209 8146 213
rect 8230 209 8264 213
rect 8321 181 8355 375
rect 8412 343 8446 347
rect 8530 343 8564 347
rect 8406 331 8452 343
rect 8406 225 8412 331
rect 8446 225 8452 331
rect 8406 213 8452 225
rect 8524 331 8570 343
rect 8524 225 8530 331
rect 8564 225 8570 331
rect 8524 213 8570 225
rect 8412 209 8446 213
rect 8530 209 8564 213
rect 8621 181 8655 375
rect 8712 343 8746 347
rect 8830 343 8864 347
rect 8706 331 8752 343
rect 8706 225 8712 331
rect 8746 225 8752 331
rect 8706 213 8752 225
rect 8824 331 8870 343
rect 8824 225 8830 331
rect 8864 225 8870 331
rect 8824 213 8870 225
rect 8712 209 8746 213
rect 8830 209 8864 213
rect 8921 181 8955 375
rect 9012 343 9046 347
rect 9130 343 9164 347
rect 9006 331 9052 343
rect 9006 225 9012 331
rect 9046 225 9052 331
rect 9006 213 9052 225
rect 9124 331 9170 343
rect 9124 225 9130 331
rect 9164 225 9170 331
rect 9124 213 9170 225
rect 9012 209 9046 213
rect 9130 209 9164 213
rect 9221 181 9255 375
rect 9312 343 9346 347
rect 9430 343 9464 347
rect 9306 331 9352 343
rect 9306 225 9312 331
rect 9346 225 9352 331
rect 9306 213 9352 225
rect 9424 331 9470 343
rect 9424 225 9430 331
rect 9464 225 9470 331
rect 9424 213 9470 225
rect 9312 209 9346 213
rect 9430 209 9464 213
rect 9521 181 9555 375
rect 9612 343 9646 347
rect 9730 343 9764 347
rect 9606 331 9652 343
rect 9606 225 9612 331
rect 9646 225 9652 331
rect 9606 213 9652 225
rect 9724 331 9770 343
rect 9724 225 9730 331
rect 9764 225 9770 331
rect 9724 213 9770 225
rect 9612 209 9646 213
rect 9730 209 9764 213
rect 9821 181 9855 375
rect 9912 343 9946 347
rect 10030 343 10064 347
rect 9906 331 9952 343
rect 9906 225 9912 331
rect 9946 225 9952 331
rect 9906 213 9952 225
rect 10024 331 10070 343
rect 10024 225 10030 331
rect 10064 225 10070 331
rect 10024 213 10070 225
rect 9912 209 9946 213
rect 10030 209 10064 213
rect 10121 181 10155 375
rect 10212 343 10246 347
rect 10330 343 10364 347
rect 10206 331 10252 343
rect 10206 225 10212 331
rect 10246 225 10252 331
rect 10206 213 10252 225
rect 10324 331 10370 343
rect 10324 225 10330 331
rect 10364 225 10370 331
rect 10324 213 10370 225
rect 10212 209 10246 213
rect 10330 209 10364 213
rect 10421 181 10455 375
rect 10512 343 10546 347
rect 10630 343 10664 347
rect 10506 331 10552 343
rect 10506 225 10512 331
rect 10546 225 10552 331
rect 10506 213 10552 225
rect 10624 331 10670 343
rect 10624 225 10630 331
rect 10664 225 10670 331
rect 10624 213 10670 225
rect 10512 209 10546 213
rect 10630 209 10664 213
rect 10721 181 10755 375
rect 10812 343 10846 347
rect 10930 343 10964 347
rect 10806 331 10852 343
rect 10806 225 10812 331
rect 10846 225 10852 331
rect 10806 213 10852 225
rect 10924 331 10970 343
rect 10924 225 10930 331
rect 10964 225 10970 331
rect 10924 213 10970 225
rect 10812 209 10846 213
rect 10930 209 10964 213
rect 11021 181 11055 375
rect 11112 343 11146 347
rect 11230 343 11264 347
rect 11106 331 11152 343
rect 11106 225 11112 331
rect 11146 225 11152 331
rect 11106 213 11152 225
rect 11224 331 11270 343
rect 11224 225 11230 331
rect 11264 225 11270 331
rect 11224 213 11270 225
rect 11112 209 11146 213
rect 11230 209 11264 213
rect 11321 181 11355 375
rect 11412 343 11446 347
rect 11530 343 11564 347
rect 11406 331 11452 343
rect 11406 225 11412 331
rect 11446 225 11452 331
rect 11406 213 11452 225
rect 11524 331 11570 343
rect 11524 225 11530 331
rect 11564 225 11570 331
rect 11524 213 11570 225
rect 11412 209 11446 213
rect 11530 209 11564 213
rect 11621 181 11655 375
rect 11712 343 11746 347
rect 11830 343 11864 347
rect 11706 331 11752 343
rect 11706 225 11712 331
rect 11746 225 11752 331
rect 11706 213 11752 225
rect 11824 331 11870 343
rect 11824 225 11830 331
rect 11864 225 11870 331
rect 11824 213 11870 225
rect 11712 209 11746 213
rect 11830 209 11864 213
rect 11921 181 11955 375
rect 12012 343 12046 347
rect 12130 343 12164 347
rect 12006 331 12052 343
rect 12006 225 12012 331
rect 12046 225 12052 331
rect 12006 213 12052 225
rect 12124 331 12170 343
rect 12124 225 12130 331
rect 12164 225 12170 331
rect 12124 213 12170 225
rect 12012 209 12046 213
rect 12130 209 12164 213
rect 12221 181 12255 375
rect 12312 343 12346 347
rect 12430 343 12464 347
rect 12306 331 12352 343
rect 12306 225 12312 331
rect 12346 225 12352 331
rect 12306 213 12352 225
rect 12424 331 12470 343
rect 12424 225 12430 331
rect 12464 225 12470 331
rect 12424 213 12470 225
rect 12312 209 12346 213
rect 12430 209 12464 213
rect 12521 181 12555 375
rect 12612 343 12646 347
rect 12730 343 12764 347
rect 12606 331 12652 343
rect 12606 225 12612 331
rect 12646 225 12652 331
rect 12606 213 12652 225
rect 12724 331 12770 343
rect 12724 225 12730 331
rect 12764 225 12770 331
rect 12724 213 12770 225
rect 12612 209 12646 213
rect 12730 209 12764 213
rect 12821 181 12855 375
rect 12912 343 12946 347
rect 13030 343 13064 347
rect 12906 331 12952 343
rect 12906 225 12912 331
rect 12946 225 12952 331
rect 12906 213 12952 225
rect 13024 331 13070 343
rect 13024 225 13030 331
rect 13064 225 13070 331
rect 13024 213 13070 225
rect 12912 209 12946 213
rect 13030 209 13064 213
rect 13121 181 13155 375
rect 13212 343 13246 347
rect 13330 343 13364 347
rect 13206 331 13252 343
rect 13206 225 13212 331
rect 13246 225 13252 331
rect 13206 213 13252 225
rect 13324 331 13370 343
rect 13324 225 13330 331
rect 13364 225 13370 331
rect 13324 213 13370 225
rect 13212 209 13246 213
rect 13330 209 13364 213
rect 13421 181 13455 375
rect 13512 343 13546 347
rect 13630 343 13664 347
rect 13506 331 13552 343
rect 13506 225 13512 331
rect 13546 225 13552 331
rect 13506 213 13552 225
rect 13624 331 13670 343
rect 13624 225 13630 331
rect 13664 225 13670 331
rect 13624 213 13670 225
rect 13512 209 13546 213
rect 13630 209 13664 213
rect 13721 181 13755 375
rect 13812 343 13846 347
rect 13930 343 13964 347
rect 13806 331 13852 343
rect 13806 225 13812 331
rect 13846 225 13852 331
rect 13806 213 13852 225
rect 13924 331 13970 343
rect 13924 225 13930 331
rect 13964 225 13970 331
rect 13924 213 13970 225
rect 13812 209 13846 213
rect 13930 209 13964 213
rect 14021 181 14055 375
rect 14112 343 14146 347
rect 14230 343 14264 347
rect 14106 331 14152 343
rect 14106 225 14112 331
rect 14146 225 14152 331
rect 14106 213 14152 225
rect 14224 331 14270 343
rect 14224 225 14230 331
rect 14264 225 14270 331
rect 14224 213 14270 225
rect 14112 209 14146 213
rect 14230 209 14264 213
rect 14321 181 14355 375
rect 14412 343 14446 347
rect 14530 343 14564 347
rect 14406 331 14452 343
rect 14406 225 14412 331
rect 14446 225 14452 331
rect 14406 213 14452 225
rect 14524 331 14570 343
rect 14524 225 14530 331
rect 14564 225 14570 331
rect 14524 213 14570 225
rect 14412 209 14446 213
rect 14530 209 14564 213
rect 14621 181 14655 375
rect 14712 343 14746 347
rect 14830 343 14864 347
rect 14706 331 14752 343
rect 14706 225 14712 331
rect 14746 225 14752 331
rect 14706 213 14752 225
rect 14824 331 14870 343
rect 14824 225 14830 331
rect 14864 225 14870 331
rect 14824 213 14870 225
rect 14712 209 14746 213
rect 14830 209 14864 213
rect 14921 181 14955 375
rect 15012 343 15046 347
rect 15130 343 15164 347
rect 15006 331 15052 343
rect 15006 225 15012 331
rect 15046 225 15052 331
rect 15006 213 15052 225
rect 15124 331 15170 343
rect 15124 225 15130 331
rect 15164 225 15170 331
rect 15124 213 15170 225
rect 15012 209 15046 213
rect 15130 209 15164 213
rect 15221 181 15255 375
rect 15312 343 15346 347
rect 15306 331 15352 343
rect 15306 225 15312 331
rect 15346 225 15352 331
rect 15306 213 15352 225
rect 15312 209 15346 213
rect 192 175 284 181
rect 192 141 204 175
rect 272 141 284 175
rect 192 135 284 141
rect 492 175 584 181
rect 492 141 504 175
rect 572 141 584 175
rect 492 135 584 141
rect 792 175 884 181
rect 792 141 804 175
rect 872 141 884 175
rect 792 135 884 141
rect 1092 175 1184 181
rect 1092 141 1104 175
rect 1172 141 1184 175
rect 1092 135 1184 141
rect 1392 175 1484 181
rect 1392 141 1404 175
rect 1472 141 1484 175
rect 1392 135 1484 141
rect 1692 175 1784 181
rect 1692 141 1704 175
rect 1772 141 1784 175
rect 1692 135 1784 141
rect 1992 175 2084 181
rect 1992 141 2004 175
rect 2072 141 2084 175
rect 1992 135 2084 141
rect 2292 175 2384 181
rect 2292 141 2304 175
rect 2372 141 2384 175
rect 2292 135 2384 141
rect 2592 175 2684 181
rect 2592 141 2604 175
rect 2672 141 2684 175
rect 2592 135 2684 141
rect 2892 175 2984 181
rect 2892 141 2904 175
rect 2972 141 2984 175
rect 2892 135 2984 141
rect 3192 175 3284 181
rect 3192 141 3204 175
rect 3272 141 3284 175
rect 3192 135 3284 141
rect 3492 175 3584 181
rect 3492 141 3504 175
rect 3572 141 3584 175
rect 3492 135 3584 141
rect 3792 175 3884 181
rect 3792 141 3804 175
rect 3872 141 3884 175
rect 3792 135 3884 141
rect 4092 175 4184 181
rect 4092 141 4104 175
rect 4172 141 4184 175
rect 4092 135 4184 141
rect 4392 175 4484 181
rect 4392 141 4404 175
rect 4472 141 4484 175
rect 4392 135 4484 141
rect 4692 175 4784 181
rect 4692 141 4704 175
rect 4772 141 4784 175
rect 4692 135 4784 141
rect 4992 175 5084 181
rect 4992 141 5004 175
rect 5072 141 5084 175
rect 4992 135 5084 141
rect 5292 175 5384 181
rect 5292 141 5304 175
rect 5372 141 5384 175
rect 5292 135 5384 141
rect 5592 175 5684 181
rect 5592 141 5604 175
rect 5672 141 5684 175
rect 5592 135 5684 141
rect 5892 175 5984 181
rect 5892 141 5904 175
rect 5972 141 5984 175
rect 5892 135 5984 141
rect 6192 175 6284 181
rect 6192 141 6204 175
rect 6272 141 6284 175
rect 6192 135 6284 141
rect 6492 175 6584 181
rect 6492 141 6504 175
rect 6572 141 6584 175
rect 6492 135 6584 141
rect 6792 175 6884 181
rect 6792 141 6804 175
rect 6872 141 6884 175
rect 6792 135 6884 141
rect 7092 175 7184 181
rect 7092 141 7104 175
rect 7172 141 7184 175
rect 7092 135 7184 141
rect 7392 175 7484 181
rect 7392 141 7404 175
rect 7472 141 7484 175
rect 7392 135 7484 141
rect 7692 175 7784 181
rect 7692 141 7704 175
rect 7772 141 7784 175
rect 7692 135 7784 141
rect 7992 175 8084 181
rect 7992 141 8004 175
rect 8072 141 8084 175
rect 7992 135 8084 141
rect 8292 175 8384 181
rect 8292 141 8304 175
rect 8372 141 8384 175
rect 8292 135 8384 141
rect 8592 175 8684 181
rect 8592 141 8604 175
rect 8672 141 8684 175
rect 8592 135 8684 141
rect 8892 175 8984 181
rect 8892 141 8904 175
rect 8972 141 8984 175
rect 8892 135 8984 141
rect 9192 175 9284 181
rect 9192 141 9204 175
rect 9272 141 9284 175
rect 9192 135 9284 141
rect 9492 175 9584 181
rect 9492 141 9504 175
rect 9572 141 9584 175
rect 9492 135 9584 141
rect 9792 175 9884 181
rect 9792 141 9804 175
rect 9872 141 9884 175
rect 9792 135 9884 141
rect 10092 175 10184 181
rect 10092 141 10104 175
rect 10172 141 10184 175
rect 10092 135 10184 141
rect 10392 175 10484 181
rect 10392 141 10404 175
rect 10472 141 10484 175
rect 10392 135 10484 141
rect 10692 175 10784 181
rect 10692 141 10704 175
rect 10772 141 10784 175
rect 10692 135 10784 141
rect 10992 175 11084 181
rect 10992 141 11004 175
rect 11072 141 11084 175
rect 10992 135 11084 141
rect 11292 175 11384 181
rect 11292 141 11304 175
rect 11372 141 11384 175
rect 11292 135 11384 141
rect 11592 175 11684 181
rect 11592 141 11604 175
rect 11672 141 11684 175
rect 11592 135 11684 141
rect 11892 175 11984 181
rect 11892 141 11904 175
rect 11972 141 11984 175
rect 11892 135 11984 141
rect 12192 175 12284 181
rect 12192 141 12204 175
rect 12272 141 12284 175
rect 12192 135 12284 141
rect 12492 175 12584 181
rect 12492 141 12504 175
rect 12572 141 12584 175
rect 12492 135 12584 141
rect 12792 175 12884 181
rect 12792 141 12804 175
rect 12872 141 12884 175
rect 12792 135 12884 141
rect 13092 175 13184 181
rect 13092 141 13104 175
rect 13172 141 13184 175
rect 13092 135 13184 141
rect 13392 175 13484 181
rect 13392 141 13404 175
rect 13472 141 13484 175
rect 13392 135 13484 141
rect 13692 175 13784 181
rect 13692 141 13704 175
rect 13772 141 13784 175
rect 13692 135 13784 141
rect 13992 175 14084 181
rect 13992 141 14004 175
rect 14072 141 14084 175
rect 13992 135 14084 141
rect 14292 175 14384 181
rect 14292 141 14304 175
rect 14372 141 14384 175
rect 14292 135 14384 141
rect 14592 175 14684 181
rect 14592 141 14604 175
rect 14672 141 14684 175
rect 14592 135 14684 141
rect 14892 175 14984 181
rect 14892 141 14904 175
rect 14972 141 14984 175
rect 14892 135 14984 141
rect 15192 175 15284 181
rect 15192 141 15204 175
rect 15272 141 15284 175
rect 15192 135 15284 141
rect 88 82 15388 94
rect 88 48 124 82
rect 352 48 424 82
rect 652 48 724 82
rect 952 48 1024 82
rect 1252 48 1324 82
rect 1552 48 1624 82
rect 1852 48 1924 82
rect 2152 48 2224 82
rect 2452 48 2524 82
rect 2752 48 2824 82
rect 3052 48 3124 82
rect 3352 48 3424 82
rect 3652 48 3724 82
rect 3952 48 4024 82
rect 4252 48 4324 82
rect 4552 48 4624 82
rect 4852 48 4924 82
rect 5152 48 5224 82
rect 5452 48 5524 82
rect 5752 48 5824 82
rect 6052 48 6124 82
rect 6352 48 6424 82
rect 6652 48 6724 82
rect 6952 48 7024 82
rect 7252 48 7324 82
rect 7552 48 7624 82
rect 7852 48 7924 82
rect 8152 48 8224 82
rect 8452 48 8524 82
rect 8752 48 8824 82
rect 9052 48 9124 82
rect 9352 48 9424 82
rect 9652 48 9724 82
rect 9952 48 10024 82
rect 10252 48 10324 82
rect 10552 48 10624 82
rect 10852 48 10924 82
rect 11152 48 11224 82
rect 11452 48 11524 82
rect 11752 48 11824 82
rect 12052 48 12124 82
rect 12352 48 12424 82
rect 12652 48 12724 82
rect 12952 48 13024 82
rect 13252 48 13324 82
rect 13552 48 13624 82
rect 13852 48 13924 82
rect 14152 48 14224 82
rect 14452 48 14524 82
rect 14752 48 14824 82
rect 15052 48 15124 82
rect 15352 48 15388 82
rect 88 36 15388 48
<< labels >>
flabel metal1 88 1168 15388 1226 0 FreeSans 256 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal1 88 36 15388 94 0 FreeSans 256 0 0 0 VSS
port 1 nsew ground bidirectional
<< end >>
