magic
tech sky130A
magscale 1 2
timestamp 1748333780
<< locali >>
rect 150 7238 250 7250
rect 150 6646 156 7238
rect 244 6646 250 7238
rect 150 6634 250 6646
rect 5572 7238 5672 7250
rect 5572 6646 5578 7238
rect 5666 6646 5672 7238
rect 5572 6634 5672 6646
rect 150 6254 253 6266
rect 150 5414 156 6254
rect 244 5414 253 6254
rect 150 5402 253 5414
rect 5572 6254 5672 6266
rect 5572 5414 5578 6254
rect 5666 5414 5672 6254
rect 5572 5402 5672 5414
rect 0 5022 112 5034
rect 0 2372 6 5022
rect 106 2372 112 5022
rect 0 2360 112 2372
rect 5710 5022 5822 5034
rect 5710 2372 5716 5022
rect 5816 2372 5822 5022
rect 5710 2360 5822 2372
rect 150 1980 253 1992
rect 150 1140 156 1980
rect 244 1140 253 1980
rect 150 1128 253 1140
rect 5572 1980 5672 1992
rect 5572 1140 5578 1980
rect 5666 1140 5672 1980
rect 5572 1128 5672 1140
rect 150 748 250 760
rect 150 156 156 748
rect 244 156 250 748
rect 150 144 250 156
rect 5572 748 5672 760
rect 5572 156 5578 748
rect 5666 156 5672 748
rect 5572 144 5672 156
<< viali >>
rect 156 6646 244 7238
rect 5578 6646 5666 7238
rect 156 5414 244 6254
rect 5578 5414 5666 6254
rect 6 2372 106 5022
rect 5716 2372 5816 5022
rect 156 1140 244 1980
rect 5578 1140 5666 1980
rect 156 156 244 748
rect 5578 156 5666 748
<< metal1 >>
rect 0 7238 250 7250
rect 0 6646 6 7238
rect 94 6646 156 7238
rect 244 6646 250 7238
rect 0 6634 250 6646
rect 5572 7238 5822 7250
rect 5572 6646 5578 7238
rect 5666 6646 5728 7238
rect 5816 6646 5822 7238
rect 5572 6634 5822 6646
rect 150 6254 250 6266
rect 150 5414 156 6254
rect 244 5414 250 6254
rect 150 5402 250 5414
rect 5572 6254 5672 6266
rect 5572 5414 5578 6254
rect 5666 5414 5672 6254
rect 5572 5402 5672 5414
rect 0 5022 112 5034
rect 0 2372 6 5022
rect 106 4988 112 5022
rect 5710 5022 5822 5034
rect 5710 4988 5716 5022
rect 106 4807 456 4988
rect 106 4737 386 4807
rect 106 4556 456 4737
rect 552 4807 788 4988
rect 552 4737 635 4807
rect 705 4737 788 4807
rect 552 4556 788 4737
rect 884 4807 1120 4988
rect 884 4737 967 4807
rect 1037 4737 1120 4807
rect 884 4556 1120 4737
rect 1216 4807 1452 4988
rect 1216 4737 1299 4807
rect 1369 4737 1452 4807
rect 1216 4556 1452 4737
rect 1548 4807 1784 4988
rect 1548 4737 1631 4807
rect 1701 4737 1784 4807
rect 1548 4556 1784 4737
rect 1880 4807 2116 4988
rect 1880 4737 1963 4807
rect 2033 4737 2116 4807
rect 1880 4556 2116 4737
rect 2212 4807 2448 4988
rect 2212 4737 2295 4807
rect 2365 4737 2448 4807
rect 2212 4556 2448 4737
rect 2544 4807 2780 4988
rect 2544 4737 2627 4807
rect 2697 4737 2780 4807
rect 2544 4556 2780 4737
rect 106 2838 112 4556
rect 2876 3472 2946 4988
rect 3042 4512 3112 4988
rect 3208 4807 3444 4988
rect 3208 4737 3291 4807
rect 3361 4737 3444 4807
rect 3208 4556 3444 4737
rect 3540 4807 3776 4988
rect 3540 4737 3623 4807
rect 3693 4737 3776 4807
rect 3540 4556 3776 4737
rect 3872 4807 4108 4988
rect 3872 4737 3955 4807
rect 4025 4737 4108 4807
rect 3872 4556 4108 4737
rect 4204 4807 4440 4988
rect 4204 4737 4287 4807
rect 4357 4737 4440 4807
rect 4204 4556 4440 4737
rect 4536 4807 4772 4988
rect 4536 4737 4619 4807
rect 4689 4737 4772 4807
rect 4536 4556 4772 4737
rect 4868 4807 5104 4988
rect 4868 4737 4951 4807
rect 5021 4737 5104 4807
rect 4868 4556 5104 4737
rect 5200 4807 5436 4988
rect 5200 4737 5283 4807
rect 5353 4737 5436 4807
rect 5200 4556 5436 4737
rect 5532 4556 5716 4988
rect 3042 4436 3112 4442
rect 2870 3402 2876 3472
rect 2946 3402 2952 3472
rect 5710 2838 5716 4556
rect 106 2406 290 2838
rect 386 2657 622 2838
rect 386 2587 469 2657
rect 539 2587 622 2657
rect 386 2406 622 2587
rect 718 2657 954 2838
rect 718 2587 801 2657
rect 871 2587 954 2657
rect 718 2406 954 2587
rect 1050 2657 1286 2838
rect 1050 2587 1133 2657
rect 1203 2587 1286 2657
rect 1050 2406 1286 2587
rect 1382 2657 1618 2838
rect 1382 2587 1465 2657
rect 1535 2587 1618 2657
rect 1382 2406 1618 2587
rect 1714 2657 1950 2838
rect 1714 2587 1797 2657
rect 1867 2587 1950 2657
rect 1714 2406 1950 2587
rect 2046 2657 2282 2838
rect 2046 2587 2129 2657
rect 2199 2587 2282 2657
rect 2046 2406 2282 2587
rect 2378 2657 2614 2838
rect 2378 2587 2461 2657
rect 2531 2587 2614 2657
rect 2378 2406 2614 2587
rect 2710 2657 2946 2838
rect 2710 2587 2793 2657
rect 2863 2587 2946 2657
rect 2710 2406 2946 2587
rect 3042 2657 3278 2838
rect 3042 2587 3125 2657
rect 3195 2587 3278 2657
rect 3042 2406 3278 2587
rect 3374 2657 3610 2838
rect 3374 2587 3457 2657
rect 3527 2587 3610 2657
rect 3374 2406 3610 2587
rect 3706 2657 3942 2838
rect 3706 2587 3789 2657
rect 3859 2587 3942 2657
rect 3706 2406 3942 2587
rect 4038 2657 4274 2838
rect 4038 2587 4121 2657
rect 4191 2587 4274 2657
rect 4038 2406 4274 2587
rect 4370 2657 4606 2838
rect 4370 2587 4453 2657
rect 4523 2587 4606 2657
rect 4370 2406 4606 2587
rect 4702 2657 4938 2838
rect 4702 2587 4785 2657
rect 4855 2587 4938 2657
rect 4702 2406 4938 2587
rect 5034 2657 5270 2838
rect 5034 2587 5117 2657
rect 5187 2587 5270 2657
rect 5034 2406 5270 2587
rect 5366 2657 5436 2838
rect 5366 2406 5436 2587
rect 5532 2406 5716 2838
rect 106 2372 112 2406
rect 0 2360 112 2372
rect 5710 2372 5716 2406
rect 5816 2372 5822 5022
rect 5710 2360 5822 2372
rect 150 1980 250 1992
rect 150 1140 156 1980
rect 244 1140 250 1980
rect 150 1128 250 1140
rect 5572 1980 5672 1992
rect 5572 1140 5578 1980
rect 5666 1140 5672 1980
rect 5572 1128 5672 1140
rect 0 748 250 760
rect 0 156 6 748
rect 94 156 156 748
rect 244 156 250 748
rect 0 144 250 156
rect 5572 748 5822 760
rect 5572 156 5578 748
rect 5666 156 5728 748
rect 5816 156 5822 748
rect 5572 144 5822 156
<< via1 >>
rect 6 6646 94 7238
rect 5728 6646 5816 7238
rect 156 5414 244 6254
rect 5578 5414 5666 6254
rect 6 2372 94 5022
rect 386 4737 456 4807
rect 635 4737 705 4807
rect 967 4737 1037 4807
rect 1299 4737 1369 4807
rect 1631 4737 1701 4807
rect 1963 4737 2033 4807
rect 2295 4737 2365 4807
rect 2627 4737 2697 4807
rect 3291 4737 3361 4807
rect 3623 4737 3693 4807
rect 3955 4737 4025 4807
rect 4287 4737 4357 4807
rect 4619 4737 4689 4807
rect 4951 4737 5021 4807
rect 5283 4737 5353 4807
rect 3042 4442 3112 4512
rect 2876 3402 2946 3472
rect 469 2587 539 2657
rect 801 2587 871 2657
rect 1133 2587 1203 2657
rect 1465 2587 1535 2657
rect 1797 2587 1867 2657
rect 2129 2587 2199 2657
rect 2461 2587 2531 2657
rect 2793 2587 2863 2657
rect 3125 2587 3195 2657
rect 3457 2587 3527 2657
rect 3789 2587 3859 2657
rect 4121 2587 4191 2657
rect 4453 2587 4523 2657
rect 4785 2587 4855 2657
rect 5117 2587 5187 2657
rect 5366 2587 5436 2657
rect 5728 2372 5816 5022
rect 156 1140 244 1980
rect 5578 1140 5666 1980
rect 6 156 94 748
rect 5728 156 5816 748
<< metal2 >>
rect 0 7238 100 7394
rect 0 6646 6 7238
rect 94 6646 100 7238
rect 0 5022 100 6646
rect 0 2372 6 5022
rect 94 2372 100 5022
rect 0 748 100 2372
rect 0 156 6 748
rect 94 156 100 748
rect 0 0 100 156
rect 150 6254 250 7394
rect 685 6709 823 7352
rect 961 6881 1099 7019
rect 1237 6881 1375 7019
rect 1513 6881 1651 7019
rect 1789 6881 1927 7019
rect 2065 6881 2203 7019
rect 2341 6881 2479 7019
rect 2617 6881 2755 7019
rect 2893 6881 3031 7019
rect 3169 6881 3307 7019
rect 3445 6881 3583 7019
rect 3721 6881 3859 7019
rect 3997 6881 4135 7019
rect 4273 6881 4411 7019
rect 4549 6881 4687 7019
rect 4825 6881 4963 7019
rect 5101 6881 5239 7019
rect 961 6837 1099 6847
rect 961 6719 971 6837
rect 1089 6719 1099 6837
rect 961 6709 1099 6719
rect 1237 6837 1375 6847
rect 1237 6719 1247 6837
rect 1365 6719 1375 6837
rect 1237 6709 1375 6719
rect 1513 6837 1651 6847
rect 1513 6719 1523 6837
rect 1641 6719 1651 6837
rect 1513 6709 1651 6719
rect 1789 6837 1927 6847
rect 1789 6719 1799 6837
rect 1917 6719 1927 6837
rect 1789 6709 1927 6719
rect 2065 6837 2203 6847
rect 2065 6719 2075 6837
rect 2193 6719 2203 6837
rect 2065 6709 2203 6719
rect 2341 6837 2479 6847
rect 2341 6719 2351 6837
rect 2469 6719 2479 6837
rect 2341 6709 2479 6719
rect 2617 6837 2755 6847
rect 2617 6719 2627 6837
rect 2745 6719 2755 6837
rect 2617 6709 2755 6719
rect 2893 6837 3031 6847
rect 2893 6719 2903 6837
rect 3021 6719 3031 6837
rect 2893 6709 3031 6719
rect 3169 6837 3307 6847
rect 3169 6719 3179 6837
rect 3297 6719 3307 6837
rect 3169 6709 3307 6719
rect 3445 6837 3583 6847
rect 3445 6719 3455 6837
rect 3573 6719 3583 6837
rect 3445 6709 3583 6719
rect 3721 6837 3859 6847
rect 3721 6719 3731 6837
rect 3849 6719 3859 6837
rect 3721 6709 3859 6719
rect 3997 6837 4135 6847
rect 3997 6719 4007 6837
rect 4125 6719 4135 6837
rect 3997 6709 4135 6719
rect 4273 6837 4411 6847
rect 4273 6719 4283 6837
rect 4401 6719 4411 6837
rect 4273 6709 4411 6719
rect 4549 6837 4687 6847
rect 4549 6719 4559 6837
rect 4677 6719 4687 6837
rect 4549 6709 4687 6719
rect 4825 6837 4963 6847
rect 4825 6719 4835 6837
rect 4953 6719 4963 6837
rect 4825 6709 4963 6719
rect 5101 6837 5239 6847
rect 5101 6719 5111 6837
rect 5229 6719 5239 6837
rect 5101 6709 5239 6719
rect 150 5414 156 6254
rect 244 5414 250 6254
rect 5572 6254 5672 7394
rect 583 5703 721 6201
rect 893 6167 963 6176
rect 893 6088 963 6097
rect 1169 6167 1239 6176
rect 1169 6088 1239 6097
rect 1445 6167 1515 6176
rect 1445 6088 1515 6097
rect 1721 6167 1791 6176
rect 1721 6088 1791 6097
rect 1997 6167 2067 6176
rect 1997 6088 2067 6097
rect 2273 6167 2343 6176
rect 2273 6088 2343 6097
rect 2549 6167 2619 6176
rect 2549 6088 2619 6097
rect 2825 6167 2895 6176
rect 2825 6088 2895 6097
rect 3101 6167 3171 6176
rect 3101 6088 3171 6097
rect 3377 6167 3447 6176
rect 3377 6088 3447 6097
rect 3653 6167 3723 6176
rect 3653 6088 3723 6097
rect 3929 6167 3999 6176
rect 3929 6088 3999 6097
rect 4205 6167 4275 6176
rect 4205 6088 4275 6097
rect 4481 6167 4551 6176
rect 4481 6088 4551 6097
rect 4757 6167 4827 6176
rect 4757 6088 4827 6097
rect 5033 6167 5103 6176
rect 5033 6088 5103 6097
rect 150 3467 250 5414
rect 5572 5414 5578 6254
rect 5666 5414 5672 6254
rect 4453 5238 4523 5243
rect 4619 5238 4689 5243
rect 4785 5238 4855 5243
rect 4951 5238 5021 5243
rect 5117 5238 5187 5243
rect 5283 5238 5353 5243
rect 4449 5178 4458 5238
rect 4518 5178 4527 5238
rect 4615 5178 4624 5238
rect 4684 5178 4693 5238
rect 4781 5178 4790 5238
rect 4850 5178 4859 5238
rect 4947 5178 4956 5238
rect 5016 5178 5025 5238
rect 5113 5178 5122 5238
rect 5182 5178 5191 5238
rect 5279 5178 5288 5238
rect 5348 5178 5357 5238
rect 4287 5157 4357 5162
rect 4283 5097 4292 5157
rect 4352 5097 4361 5157
rect 4121 5027 4191 5032
rect 4117 4967 4126 5027
rect 4186 4967 4195 5027
rect 3955 4897 4025 4902
rect 3951 4837 3960 4897
rect 4020 4837 4029 4897
rect 3955 4807 4025 4837
rect 150 3407 155 3467
rect 215 3407 250 3467
rect 150 1980 250 3407
rect 303 4737 386 4807
rect 456 4737 462 4807
rect 629 4737 635 4807
rect 705 4737 711 4807
rect 961 4737 967 4807
rect 1037 4737 1043 4807
rect 1293 4737 1299 4807
rect 1369 4737 1375 4807
rect 1625 4737 1631 4807
rect 1701 4737 1707 4807
rect 1957 4737 1963 4807
rect 2033 4737 2039 4807
rect 2289 4737 2295 4807
rect 2365 4737 2371 4807
rect 2621 4737 2627 4807
rect 2697 4737 2703 4807
rect 3285 4737 3291 4807
rect 3361 4737 3367 4807
rect 3617 4737 3623 4807
rect 3693 4737 3699 4807
rect 3789 4767 3859 4772
rect 303 2216 373 4737
rect 463 2587 469 2657
rect 539 2587 545 2657
rect 469 2216 539 2587
rect 635 2216 705 4737
rect 795 2587 801 2657
rect 871 2587 877 2657
rect 801 2216 871 2587
rect 967 2216 1037 4737
rect 1127 2587 1133 2657
rect 1203 2587 1209 2657
rect 1133 2216 1203 2587
rect 1299 2216 1369 4737
rect 1459 2587 1465 2657
rect 1535 2587 1541 2657
rect 1465 2297 1535 2587
rect 1631 2427 1701 4737
rect 1963 2687 2033 4737
rect 2295 2947 2365 4737
rect 2627 3207 2697 4737
rect 2959 4442 3042 4512
rect 3112 4442 3118 4512
rect 2959 4117 3029 4442
rect 3291 4377 3361 4737
rect 3623 4637 3693 4737
rect 3785 4707 3794 4767
rect 3854 4707 3863 4767
rect 3949 4737 3955 4807
rect 4025 4737 4031 4807
rect 3619 4577 3628 4637
rect 3688 4577 3697 4637
rect 3623 4572 3693 4577
rect 3457 4507 3527 4512
rect 3453 4447 3462 4507
rect 3522 4447 3531 4507
rect 3287 4317 3296 4377
rect 3356 4317 3365 4377
rect 3291 4312 3361 4317
rect 3125 4247 3195 4252
rect 3121 4187 3130 4247
rect 3190 4187 3199 4247
rect 2955 4057 2964 4117
rect 3024 4057 3033 4117
rect 2959 3607 3029 4057
rect 2950 3537 2959 3607
rect 3029 3537 3038 3607
rect 2876 3472 2946 3478
rect 2872 3407 2876 3467
rect 2946 3407 2950 3467
rect 2876 3396 2946 3402
rect 2793 3337 2863 3342
rect 2789 3277 2798 3337
rect 2858 3277 2867 3337
rect 2623 3147 2632 3207
rect 2692 3147 2701 3207
rect 2627 3142 2697 3147
rect 2461 3077 2531 3082
rect 2457 3017 2466 3077
rect 2526 3017 2535 3077
rect 2291 2887 2300 2947
rect 2360 2887 2369 2947
rect 2295 2882 2365 2887
rect 2129 2817 2199 2822
rect 2125 2757 2134 2817
rect 2194 2757 2203 2817
rect 1791 2587 1797 2657
rect 1867 2587 1873 2657
rect 1959 2627 1968 2687
rect 2028 2627 2037 2687
rect 2129 2657 2199 2757
rect 2461 2657 2531 3017
rect 2793 2657 2863 3277
rect 3125 2657 3195 4187
rect 3457 2657 3527 4447
rect 3789 2657 3859 4707
rect 4121 2657 4191 4967
rect 4287 4807 4357 5097
rect 4281 4737 4287 4807
rect 4357 4737 4363 4807
rect 4453 2657 4523 5178
rect 4619 4807 4689 5178
rect 4613 4737 4619 4807
rect 4689 4737 4695 4807
rect 4785 2657 4855 5178
rect 4951 4807 5021 5178
rect 4945 4737 4951 4807
rect 5021 4737 5027 4807
rect 5117 2657 5187 5178
rect 5283 4807 5353 5178
rect 5277 4737 5283 4807
rect 5353 4737 5359 4807
rect 5449 2657 5519 2663
rect 1963 2622 2033 2627
rect 2123 2587 2129 2657
rect 2199 2587 2205 2657
rect 2455 2587 2461 2657
rect 2531 2587 2537 2657
rect 2787 2587 2793 2657
rect 2863 2587 2869 2657
rect 3119 2587 3125 2657
rect 3195 2587 3201 2657
rect 3451 2587 3457 2657
rect 3527 2587 3533 2657
rect 3783 2587 3789 2657
rect 3859 2587 3865 2657
rect 4115 2587 4121 2657
rect 4191 2587 4197 2657
rect 4447 2587 4453 2657
rect 4523 2587 4529 2657
rect 4779 2587 4785 2657
rect 4855 2587 4861 2657
rect 5111 2587 5117 2657
rect 5187 2587 5193 2657
rect 5360 2587 5366 2657
rect 5436 2652 5519 2657
rect 5436 2592 5454 2652
rect 5514 2592 5523 2652
rect 5436 2587 5519 2592
rect 1797 2557 1867 2587
rect 5449 2581 5519 2587
rect 1793 2497 1802 2557
rect 1862 2497 1871 2557
rect 1797 2492 1867 2497
rect 1627 2367 1636 2427
rect 1696 2367 1705 2427
rect 1631 2362 1701 2367
rect 1461 2237 1470 2297
rect 1530 2237 1539 2297
rect 1465 2232 1535 2237
rect 299 2156 308 2216
rect 368 2156 377 2216
rect 465 2156 474 2216
rect 534 2156 543 2216
rect 631 2156 640 2216
rect 700 2156 709 2216
rect 797 2156 806 2216
rect 866 2156 875 2216
rect 963 2156 972 2216
rect 1032 2156 1041 2216
rect 1129 2156 1138 2216
rect 1198 2156 1207 2216
rect 1295 2156 1304 2216
rect 1364 2156 1373 2216
rect 303 2151 373 2156
rect 469 2151 539 2156
rect 635 2151 705 2156
rect 801 2151 871 2156
rect 967 2151 1037 2156
rect 1133 2151 1203 2156
rect 1299 2151 1369 2156
rect 150 1140 156 1980
rect 244 1140 250 1980
rect 5572 1980 5672 5414
rect 719 1297 789 1306
rect 719 1218 789 1227
rect 995 1297 1065 1306
rect 995 1218 1065 1227
rect 1271 1297 1341 1306
rect 1271 1218 1341 1227
rect 1547 1297 1617 1306
rect 1547 1218 1617 1227
rect 1823 1297 1893 1306
rect 1823 1218 1893 1227
rect 2099 1297 2169 1306
rect 2099 1218 2169 1227
rect 2375 1297 2445 1306
rect 2375 1218 2445 1227
rect 2651 1297 2721 1306
rect 2651 1218 2721 1227
rect 2927 1297 2997 1306
rect 2927 1218 2997 1227
rect 3203 1297 3273 1306
rect 3203 1218 3273 1227
rect 3479 1297 3549 1306
rect 3479 1218 3549 1227
rect 3755 1297 3825 1306
rect 3755 1218 3825 1227
rect 4031 1297 4101 1306
rect 4031 1218 4101 1227
rect 4307 1297 4377 1306
rect 4307 1218 4377 1227
rect 4583 1297 4653 1306
rect 4583 1218 4653 1227
rect 4859 1297 4929 1306
rect 4859 1218 4929 1227
rect 5135 1297 5205 1306
rect 5135 1218 5205 1227
rect 150 0 250 1140
rect 5572 1140 5578 1980
rect 5666 1140 5672 1980
rect 583 675 721 685
rect 583 557 593 675
rect 711 557 721 675
rect 583 547 721 557
rect 859 675 997 685
rect 859 557 869 675
rect 987 557 997 675
rect 859 547 997 557
rect 1135 675 1273 685
rect 1135 557 1145 675
rect 1263 557 1273 675
rect 1135 547 1273 557
rect 1411 675 1549 685
rect 1411 557 1421 675
rect 1539 557 1549 675
rect 1411 547 1549 557
rect 1687 675 1825 685
rect 1687 557 1697 675
rect 1815 557 1825 675
rect 1687 547 1825 557
rect 1963 675 2101 685
rect 1963 557 1973 675
rect 2091 557 2101 675
rect 1963 547 2101 557
rect 2239 675 2377 685
rect 2239 557 2249 675
rect 2367 557 2377 675
rect 2239 547 2377 557
rect 2515 675 2653 685
rect 2515 557 2525 675
rect 2643 557 2653 675
rect 2515 547 2653 557
rect 2791 675 2929 685
rect 2791 557 2801 675
rect 2919 557 2929 675
rect 2791 547 2929 557
rect 3067 675 3205 685
rect 3067 557 3077 675
rect 3195 557 3205 675
rect 3067 547 3205 557
rect 3343 675 3481 685
rect 3343 557 3353 675
rect 3471 557 3481 675
rect 3343 547 3481 557
rect 3619 675 3757 685
rect 3619 557 3629 675
rect 3747 557 3757 675
rect 3619 547 3757 557
rect 3895 675 4033 685
rect 3895 557 3905 675
rect 4023 557 4033 675
rect 3895 547 4033 557
rect 4171 675 4309 685
rect 4171 557 4181 675
rect 4299 557 4309 675
rect 4171 547 4309 557
rect 4447 675 4585 685
rect 4447 557 4457 675
rect 4575 557 4585 675
rect 4447 547 4585 557
rect 4723 675 4861 685
rect 4723 557 4733 675
rect 4851 557 4861 675
rect 4723 547 4861 557
rect 4999 675 5137 685
rect 4999 557 5009 675
rect 5127 557 5137 675
rect 4999 547 5137 557
rect 583 375 721 513
rect 859 375 997 513
rect 1135 375 1273 513
rect 1411 375 1549 513
rect 1687 375 1825 513
rect 1963 375 2101 513
rect 2239 375 2377 513
rect 2515 375 2653 513
rect 2791 375 2929 513
rect 3067 375 3205 513
rect 3343 375 3481 513
rect 3619 375 3757 513
rect 3895 375 4033 513
rect 4171 375 4309 513
rect 4447 375 4585 513
rect 4723 375 4861 513
rect 4999 375 5137 513
rect 5572 0 5672 1140
rect 5722 7238 5822 7394
rect 5722 6646 5728 7238
rect 5816 6646 5822 7238
rect 5722 5022 5822 6646
rect 5722 2372 5728 5022
rect 5816 2372 5822 5022
rect 5722 748 5822 2372
rect 5722 156 5728 748
rect 5816 156 5822 748
rect 5722 0 5822 156
<< via2 >>
rect 971 6719 1089 6837
rect 1247 6719 1365 6837
rect 1523 6719 1641 6837
rect 1799 6719 1917 6837
rect 2075 6719 2193 6837
rect 2351 6719 2469 6837
rect 2627 6719 2745 6837
rect 2903 6719 3021 6837
rect 3179 6719 3297 6837
rect 3455 6719 3573 6837
rect 3731 6719 3849 6837
rect 4007 6719 4125 6837
rect 4283 6719 4401 6837
rect 4559 6719 4677 6837
rect 4835 6719 4953 6837
rect 5111 6719 5229 6837
rect 893 6097 963 6167
rect 1169 6097 1239 6167
rect 1445 6097 1515 6167
rect 1721 6097 1791 6167
rect 1997 6097 2067 6167
rect 2273 6097 2343 6167
rect 2549 6097 2619 6167
rect 2825 6097 2895 6167
rect 3101 6097 3171 6167
rect 3377 6097 3447 6167
rect 3653 6097 3723 6167
rect 3929 6097 3999 6167
rect 4205 6097 4275 6167
rect 4481 6097 4551 6167
rect 4757 6097 4827 6167
rect 5033 6097 5103 6167
rect 4458 5178 4518 5238
rect 4624 5178 4684 5238
rect 4790 5178 4850 5238
rect 4956 5178 5016 5238
rect 5122 5178 5182 5238
rect 5288 5178 5348 5238
rect 4292 5097 4352 5157
rect 4126 4967 4186 5027
rect 3960 4837 4020 4897
rect 155 3407 215 3467
rect 3794 4707 3854 4767
rect 3628 4577 3688 4637
rect 3462 4447 3522 4507
rect 3296 4317 3356 4377
rect 3130 4187 3190 4247
rect 2964 4057 3024 4117
rect 2959 3537 3029 3607
rect 2881 3407 2941 3467
rect 2798 3277 2858 3337
rect 2632 3147 2692 3207
rect 2466 3017 2526 3077
rect 2300 2887 2360 2947
rect 2134 2757 2194 2817
rect 1968 2627 2028 2687
rect 5454 2592 5514 2652
rect 1802 2497 1862 2557
rect 1636 2367 1696 2427
rect 1470 2237 1530 2297
rect 308 2156 368 2216
rect 474 2156 534 2216
rect 640 2156 700 2216
rect 806 2156 866 2216
rect 972 2156 1032 2216
rect 1138 2156 1198 2216
rect 1304 2156 1364 2216
rect 719 1227 789 1297
rect 995 1227 1065 1297
rect 1271 1227 1341 1297
rect 1547 1227 1617 1297
rect 1823 1227 1893 1297
rect 2099 1227 2169 1297
rect 2375 1227 2445 1297
rect 2651 1227 2721 1297
rect 2927 1227 2997 1297
rect 3203 1227 3273 1297
rect 3479 1227 3549 1297
rect 3755 1227 3825 1297
rect 4031 1227 4101 1297
rect 4307 1227 4377 1297
rect 4583 1227 4653 1297
rect 4859 1227 4929 1297
rect 5135 1227 5205 1297
rect 593 557 711 675
rect 869 557 987 675
rect 1145 557 1263 675
rect 1421 557 1539 675
rect 1697 557 1815 675
rect 1973 557 2091 675
rect 2249 557 2367 675
rect 2525 557 2643 675
rect 2801 557 2919 675
rect 3077 557 3195 675
rect 3353 557 3471 675
rect 3629 557 3747 675
rect 3905 557 4023 675
rect 4181 557 4299 675
rect 4457 557 4575 675
rect 4733 557 4851 675
rect 5009 557 5127 675
<< metal3 >>
rect 961 6837 5239 6847
rect 961 6719 971 6837
rect 1089 6719 1247 6837
rect 1365 6719 1523 6837
rect 1641 6719 1799 6837
rect 1917 6719 2075 6837
rect 2193 6719 2351 6837
rect 2469 6719 2627 6837
rect 2745 6719 2903 6837
rect 3021 6719 3179 6837
rect 3297 6719 3455 6837
rect 3573 6719 3731 6837
rect 3849 6719 4007 6837
rect 4125 6719 4283 6837
rect 4401 6719 4559 6837
rect 4677 6719 4835 6837
rect 4953 6719 5111 6837
rect 5229 6719 5239 6837
rect 961 6709 5239 6719
rect 5038 6172 5108 6178
rect 888 6167 968 6172
rect 888 6097 893 6167
rect 963 6097 968 6167
rect 888 6092 968 6097
rect 1164 6167 1244 6172
rect 1164 6097 1169 6167
rect 1239 6097 1244 6167
rect 1164 6092 1244 6097
rect 1440 6167 1520 6172
rect 1440 6097 1445 6167
rect 1515 6097 1520 6167
rect 1440 6092 1520 6097
rect 1716 6167 1796 6172
rect 1716 6097 1721 6167
rect 1791 6097 1796 6167
rect 1716 6092 1796 6097
rect 1992 6167 2072 6172
rect 1992 6097 1997 6167
rect 2067 6097 2072 6167
rect 1992 6092 2072 6097
rect 2268 6167 2348 6172
rect 2268 6097 2273 6167
rect 2343 6097 2348 6167
rect 2268 6092 2348 6097
rect 2544 6167 2624 6172
rect 2544 6097 2549 6167
rect 2619 6097 2624 6167
rect 2544 6092 2624 6097
rect 2820 6167 2900 6172
rect 2820 6097 2825 6167
rect 2895 6097 2900 6167
rect 2820 6092 2900 6097
rect 3096 6167 3176 6172
rect 3096 6097 3101 6167
rect 3171 6097 3176 6167
rect 3096 6092 3176 6097
rect 3372 6167 3452 6172
rect 3372 6097 3377 6167
rect 3447 6097 3452 6167
rect 3372 6092 3452 6097
rect 3648 6167 3728 6172
rect 3648 6097 3653 6167
rect 3723 6097 3728 6167
rect 3648 6092 3728 6097
rect 3924 6167 4004 6172
rect 3924 6097 3929 6167
rect 3999 6097 4004 6167
rect 3924 6092 4004 6097
rect 4200 6167 4280 6172
rect 4200 6097 4205 6167
rect 4275 6097 4280 6167
rect 4200 6092 4280 6097
rect 4476 6167 4556 6172
rect 4476 6097 4481 6167
rect 4551 6097 4556 6167
rect 4476 6092 4556 6097
rect 4752 6167 4832 6172
rect 4752 6097 4757 6167
rect 4827 6097 4832 6167
rect 4752 6092 4832 6097
rect 5028 6167 5108 6172
rect 5028 6097 5033 6167
rect 5103 6097 5108 6167
rect 5028 6092 5108 6097
rect 893 4122 963 6092
rect 1169 4252 1239 6092
rect 1445 4382 1515 6092
rect 1721 4512 1791 6092
rect 1997 4642 2067 6092
rect 2273 4772 2343 6092
rect 2549 4902 2619 6092
rect 2825 5032 2895 6092
rect 3101 5162 3171 6092
rect 3377 5292 3447 6092
rect 3653 5422 3723 6092
rect 3929 5552 3999 6092
rect 4205 5682 4275 6092
rect 4481 5812 4551 6092
rect 4757 5942 4827 6092
rect 5033 6077 5108 6092
rect 5033 6007 5519 6077
rect 4757 5872 5353 5942
rect 4481 5742 5187 5812
rect 4205 5612 5021 5682
rect 3929 5482 4855 5552
rect 3653 5352 4689 5422
rect 3377 5238 4523 5292
rect 3377 5222 4458 5238
rect 4453 5178 4458 5222
rect 4518 5178 4523 5238
rect 4453 5173 4523 5178
rect 4619 5238 4689 5352
rect 4619 5178 4624 5238
rect 4684 5178 4689 5238
rect 4619 5173 4689 5178
rect 4785 5238 4855 5482
rect 4785 5178 4790 5238
rect 4850 5178 4855 5238
rect 4785 5173 4855 5178
rect 4951 5238 5021 5612
rect 4951 5178 4956 5238
rect 5016 5178 5021 5238
rect 4951 5173 5021 5178
rect 5117 5238 5187 5742
rect 5117 5178 5122 5238
rect 5182 5178 5187 5238
rect 5117 5173 5187 5178
rect 5283 5238 5353 5872
rect 5283 5178 5288 5238
rect 5348 5178 5353 5238
rect 5283 5173 5353 5178
rect 3101 5157 4357 5162
rect 3101 5097 4292 5157
rect 4352 5097 4357 5157
rect 3101 5092 4357 5097
rect 2825 5027 4191 5032
rect 2825 4967 4126 5027
rect 4186 4967 4191 5027
rect 2825 4962 4191 4967
rect 2549 4897 4025 4902
rect 2549 4837 3960 4897
rect 4020 4837 4025 4897
rect 2549 4832 4025 4837
rect 2273 4767 3859 4772
rect 2273 4707 3794 4767
rect 3854 4707 3859 4767
rect 2273 4702 3859 4707
rect 1997 4637 3693 4642
rect 1997 4577 3628 4637
rect 3688 4577 3693 4637
rect 1997 4572 3693 4577
rect 1721 4507 3527 4512
rect 1721 4447 3462 4507
rect 3522 4447 3527 4507
rect 1721 4442 3527 4447
rect 1445 4377 3361 4382
rect 1445 4317 3296 4377
rect 3356 4317 3361 4377
rect 1445 4312 3361 4317
rect 1169 4247 3195 4252
rect 1169 4187 3130 4247
rect 3190 4187 3195 4247
rect 1169 4182 3195 4187
rect 893 4117 3029 4122
rect 893 4057 2964 4117
rect 3024 4057 3029 4117
rect 893 4052 3029 4057
rect 2954 3607 3034 3612
rect 2954 3537 2959 3607
rect 3029 3537 5340 3607
rect 2954 3532 3034 3537
rect 150 3467 5205 3472
rect 150 3407 155 3467
rect 215 3407 2881 3467
rect 2941 3407 5205 3467
rect 150 3402 5205 3407
rect 2793 3337 4929 3342
rect 2793 3277 2798 3337
rect 2858 3277 4929 3337
rect 2793 3272 4929 3277
rect 2627 3207 4653 3212
rect 2627 3147 2632 3207
rect 2692 3147 4653 3207
rect 2627 3142 4653 3147
rect 2461 3077 4377 3082
rect 2461 3017 2466 3077
rect 2526 3017 4377 3077
rect 2461 3012 4377 3017
rect 2295 2947 4101 2952
rect 2295 2887 2300 2947
rect 2360 2887 4101 2947
rect 2295 2882 4101 2887
rect 2129 2817 3825 2822
rect 2129 2757 2134 2817
rect 2194 2757 3825 2817
rect 2129 2752 3825 2757
rect 1963 2687 3549 2692
rect 1963 2627 1968 2687
rect 2028 2627 3549 2687
rect 1963 2622 3549 2627
rect 1797 2557 3273 2562
rect 1797 2497 1802 2557
rect 1862 2497 3273 2557
rect 1797 2492 3273 2497
rect 1631 2427 2997 2432
rect 1631 2367 1636 2427
rect 1696 2367 2997 2427
rect 1631 2362 2997 2367
rect 1465 2297 2721 2302
rect 1465 2237 1470 2297
rect 1530 2237 2721 2297
rect 1465 2232 2721 2237
rect 303 2216 373 2221
rect 303 2156 308 2216
rect 368 2156 373 2216
rect 303 1387 373 2156
rect 469 2216 539 2221
rect 469 2156 474 2216
rect 534 2156 539 2216
rect 469 1522 539 2156
rect 635 2216 705 2221
rect 635 2156 640 2216
rect 700 2156 705 2216
rect 635 1652 705 2156
rect 801 2216 871 2221
rect 801 2156 806 2216
rect 866 2156 871 2216
rect 801 1782 871 2156
rect 967 2216 1037 2221
rect 967 2156 972 2216
rect 1032 2156 1037 2216
rect 967 1912 1037 2156
rect 1133 2216 1203 2221
rect 1133 2156 1138 2216
rect 1198 2156 1203 2216
rect 1133 2042 1203 2156
rect 1299 2216 1369 2221
rect 1299 2156 1304 2216
rect 1364 2172 1369 2216
rect 1364 2156 2445 2172
rect 1299 2102 2445 2156
rect 1133 1972 2169 2042
rect 967 1842 1893 1912
rect 801 1712 1617 1782
rect 635 1582 1341 1652
rect 469 1452 1065 1522
rect 303 1317 789 1387
rect 714 1302 789 1317
rect 995 1302 1065 1452
rect 1271 1302 1341 1582
rect 1547 1302 1617 1712
rect 1823 1302 1893 1842
rect 2099 1302 2169 1972
rect 2375 1302 2445 2102
rect 2651 1302 2721 2232
rect 2927 1302 2997 2362
rect 3203 1302 3273 2492
rect 3479 1302 3549 2622
rect 3755 1302 3825 2752
rect 4031 1302 4101 2882
rect 4307 1302 4377 3012
rect 4583 1302 4653 3142
rect 4859 1302 4929 3272
rect 5135 1302 5205 3402
rect 714 1297 794 1302
rect 714 1227 719 1297
rect 789 1227 794 1297
rect 714 1222 794 1227
rect 990 1297 1070 1302
rect 990 1227 995 1297
rect 1065 1227 1070 1297
rect 990 1222 1070 1227
rect 1266 1297 1346 1302
rect 1266 1227 1271 1297
rect 1341 1227 1346 1297
rect 1266 1222 1346 1227
rect 1542 1297 1622 1302
rect 1542 1227 1547 1297
rect 1617 1227 1622 1297
rect 1542 1222 1622 1227
rect 1818 1297 1898 1302
rect 1818 1227 1823 1297
rect 1893 1227 1898 1297
rect 1818 1222 1898 1227
rect 2094 1297 2174 1302
rect 2094 1227 2099 1297
rect 2169 1227 2174 1297
rect 2094 1222 2174 1227
rect 2370 1297 2450 1302
rect 2370 1227 2375 1297
rect 2445 1227 2450 1297
rect 2370 1222 2450 1227
rect 2646 1297 2726 1302
rect 2646 1227 2651 1297
rect 2721 1227 2726 1297
rect 2646 1222 2726 1227
rect 2922 1297 3002 1302
rect 2922 1227 2927 1297
rect 2997 1227 3002 1297
rect 2922 1222 3002 1227
rect 3198 1297 3278 1302
rect 3198 1227 3203 1297
rect 3273 1227 3278 1297
rect 3198 1222 3278 1227
rect 3474 1297 3554 1302
rect 3474 1227 3479 1297
rect 3549 1227 3554 1297
rect 3474 1222 3554 1227
rect 3750 1297 3830 1302
rect 3750 1227 3755 1297
rect 3825 1227 3830 1297
rect 3750 1222 3830 1227
rect 4026 1297 4106 1302
rect 4026 1227 4031 1297
rect 4101 1227 4106 1297
rect 4026 1222 4106 1227
rect 4302 1297 4382 1302
rect 4302 1227 4307 1297
rect 4377 1227 4382 1297
rect 4302 1222 4382 1227
rect 4578 1297 4658 1302
rect 4578 1227 4583 1297
rect 4653 1227 4658 1297
rect 4578 1222 4658 1227
rect 4854 1297 4934 1302
rect 4854 1227 4859 1297
rect 4929 1227 4934 1297
rect 4854 1222 4934 1227
rect 5130 1297 5210 1302
rect 5130 1227 5135 1297
rect 5205 1227 5210 1297
rect 5130 1222 5210 1227
rect 5270 815 5340 3537
rect 5449 2662 5519 6007
rect 5444 2652 5524 2662
rect 5444 2592 5454 2652
rect 5514 2592 5524 2652
rect 5444 2582 5524 2592
rect 893 745 5340 815
rect 893 685 963 745
rect 1445 685 1515 745
rect 1997 685 2067 745
rect 2549 685 2619 745
rect 3101 685 3171 745
rect 3653 685 3723 745
rect 4205 685 4275 745
rect 4757 685 4827 745
rect 583 675 721 685
rect 583 557 593 675
rect 711 557 721 675
rect 583 547 721 557
rect 859 675 997 685
rect 859 557 869 675
rect 987 557 997 675
rect 859 547 997 557
rect 1135 675 1273 685
rect 1135 557 1145 675
rect 1263 557 1273 675
rect 1135 547 1273 557
rect 1411 675 1549 685
rect 1411 557 1421 675
rect 1539 557 1549 675
rect 1411 547 1549 557
rect 1687 675 1825 685
rect 1687 557 1697 675
rect 1815 557 1825 675
rect 1687 547 1825 557
rect 1963 675 2101 685
rect 1963 557 1973 675
rect 2091 557 2101 675
rect 1963 547 2101 557
rect 2239 675 2377 685
rect 2239 557 2249 675
rect 2367 557 2377 675
rect 2239 547 2377 557
rect 2515 675 2653 685
rect 2515 557 2525 675
rect 2643 557 2653 675
rect 2515 547 2653 557
rect 2791 675 2929 685
rect 2791 557 2801 675
rect 2919 557 2929 675
rect 2791 547 2929 557
rect 3067 675 3205 685
rect 3067 557 3077 675
rect 3195 557 3205 675
rect 3067 547 3205 557
rect 3343 675 3481 685
rect 3343 557 3353 675
rect 3471 557 3481 675
rect 3343 547 3481 557
rect 3619 675 3757 685
rect 3619 557 3629 675
rect 3747 557 3757 675
rect 3619 547 3757 557
rect 3895 675 4033 685
rect 3895 557 3905 675
rect 4023 557 4033 675
rect 3895 547 4033 557
rect 4171 675 4309 685
rect 4171 557 4181 675
rect 4299 557 4309 675
rect 4171 547 4309 557
rect 4447 675 4585 685
rect 4447 557 4457 675
rect 4575 557 4585 675
rect 4447 547 4585 557
rect 4723 675 4861 685
rect 4723 557 4733 675
rect 4851 557 4861 675
rect 4723 547 4861 557
rect 4999 675 5137 685
rect 4999 557 5009 675
rect 5127 557 5137 675
rect 4999 547 5137 557
rect 617 487 687 547
rect 1169 487 1239 547
rect 1721 487 1791 547
rect 2273 487 2343 547
rect 2825 487 2895 547
rect 3377 487 3447 547
rect 3929 487 3999 547
rect 4481 487 4551 547
rect 5033 487 5103 547
rect 5449 487 5519 2582
rect 617 417 5519 487
use passgates  passgates_0
timestamp 1748309517
transform -1 0 5681 0 -1 7394
box 0 0 5540 2076
use passgates  passgates_2
timestamp 1748309517
transform 1 0 141 0 1 0
box 0 0 5540 2076
use sky130_fd_pr__res_xhigh_po_0p35_7C4M5Y  sky130_fd_pr__res_xhigh_po_0p35_7C4M5Y_0
timestamp 1748333645
transform 1 0 2911 0 1 3697
box -2911 -1511 2911 1511
<< labels >>
flabel metal2 0 0 100 7214 1 FreeSans 400 0 0 0 VSS
port 1 n ground bidirectional
flabel metal2 150 0 250 7214 1 FreeSans 400 0 0 0 VDD
port 2 n power bidirectional
flabel metal3 617 417 5519 487 1 FreeSans 400 0 0 0 A
flabel metal3 893 745 5340 815 1 FreeSans 400 0 0 0 B
flabel metal2 583 375 721 513 1 FreeSans 400 0 0 0 C[0]
port 20 n signal default
flabel metal2 859 375 997 513 1 FreeSans 400 0 0 0 C[1]
port 21 n signal default
flabel metal2 1135 375 1273 513 1 FreeSans 400 0 0 0 C[2]
port 22 n signal default
flabel metal2 1411 375 1549 513 1 FreeSans 400 0 0 0 C[3]
port 23 n signal default
flabel metal2 1687 375 1825 513 1 FreeSans 400 0 0 0 C[4]
port 24 n signal default
flabel metal2 1963 375 2101 513 1 FreeSans 400 0 0 0 C[5]
port 25 n signal default
flabel metal2 2239 375 2377 513 1 FreeSans 400 0 0 0 C[6]
port 26 n signal default
flabel metal2 2515 375 2653 513 1 FreeSans 400 0 0 0 C[7]
port 27 n signal default
flabel metal2 2791 375 2929 513 1 FreeSans 400 0 0 0 C[8]
port 28 n signal default
flabel metal2 3067 375 3205 513 1 FreeSans 400 0 0 0 C[9]
port 29 n signal default
flabel metal2 3343 375 3481 513 1 FreeSans 400 0 0 0 C[10]
port 30 n signal default
flabel metal2 3619 375 3757 513 1 FreeSans 400 0 0 0 C[11]
port 31 n signal default
flabel metal2 3895 375 4033 513 1 FreeSans 400 0 0 0 C[12]
port 32 n signal default
flabel metal2 4171 375 4309 513 1 FreeSans 400 0 0 0 C[13]
port 33 n signal default
flabel metal2 4447 375 4585 513 1 FreeSans 400 0 0 0 C[14]
port 34 n signal default
flabel metal2 4723 375 4861 513 1 FreeSans 400 0 0 0 C[15]
port 35 n signal default
flabel metal2 4999 375 5137 513 1 FreeSans 400 0 0 0 C[16]
port 36 n signal default
flabel metal3 961 6709 5239 6847 1 FreeSans 400 0 0 0 VOUT
port 3 n signal default
flabel metal2 5101 6881 5239 7019 1 FreeSans 400 0 0 0 D[0]
port 4 n signal default
flabel metal2 4825 6881 4963 7019 1 FreeSans 400 0 0 0 D[1]
port 5 n signal default
flabel metal2 4549 6881 4687 7019 1 FreeSans 400 0 0 0 D[2]
port 6 n signal default
flabel metal2 4273 6881 4411 7019 1 FreeSans 400 0 0 0 D[3]
port 7 n signal default
flabel metal2 3997 6881 4135 7019 1 FreeSans 400 0 0 0 D[4]
port 8 n signal default
flabel metal2 3721 6881 3859 7019 1 FreeSans 400 0 0 0 D[5]
port 9 n signal default
flabel metal2 3445 6881 3583 7019 1 FreeSans 400 0 0 0 D[6]
port 10 n signal default
flabel metal2 3169 6881 3307 7019 1 FreeSans 400 0 0 0 D[7]
port 11 n signal default
flabel metal2 2893 6881 3031 7019 1 FreeSans 400 0 0 0 D[8]
port 12 n signal default
flabel metal2 2617 6881 2755 7019 1 FreeSans 400 0 0 0 D[9]
port 13 n signal default
flabel metal2 2341 6881 2479 7019 1 FreeSans 400 0 0 0 D[10]
port 14 n signal default
flabel metal2 2065 6881 2203 7019 1 FreeSans 400 0 0 0 D[11]
port 15 n signal default
flabel metal2 1789 6881 1927 7019 1 FreeSans 400 0 0 0 D[12]
port 16 n signal default
flabel metal2 1513 6881 1651 7019 1 FreeSans 400 0 0 0 D[13]
port 17 n signal default
flabel metal2 1237 6881 1375 7019 1 FreeSans 400 0 0 0 D[14]
port 18 n signal default
flabel metal2 961 6881 1099 7019 1 FreeSans 400 0 0 0 D[15]
port 19 n signal default
<< end >>
