magic
tech sky130A
magscale 1 2
timestamp 1748330861
<< dnwell >>
rect 5459 12246 22267 32733
<< nwell >>
rect 5349 32527 22377 32843
rect 5349 12452 5665 32527
rect 22061 12452 22377 32527
rect 5349 12136 22377 12452
<< mvnsubdiff >>
rect 5416 32756 22310 32776
rect 5416 32722 5496 32756
rect 22230 32722 22310 32756
rect 5416 32702 22310 32722
rect 5416 32696 5490 32702
rect 5416 12283 5436 32696
rect 5470 12283 5490 32696
rect 5416 12277 5490 12283
rect 22236 32696 22310 32702
rect 22236 12283 22256 32696
rect 22290 12283 22310 32696
rect 22236 12277 22310 12283
rect 5416 12257 22310 12277
rect 5416 12223 5496 12257
rect 22230 12223 22310 12257
rect 5416 12203 22310 12223
<< mvnsubdiffcont >>
rect 5496 32722 22230 32756
rect 5436 12283 5470 32696
rect 22256 12283 22290 32696
rect 5496 12223 22230 12257
<< locali >>
rect 5436 32722 5496 32756
rect 22230 32722 22290 32756
rect 5436 32696 5470 32722
rect 5436 12257 5470 12283
rect 22256 32696 22290 32722
rect 22256 12257 22290 12283
rect 5436 12223 5496 12257
rect 22230 12223 22290 12257
use toplevel  toplevel_0
timestamp 1748326618
transform 1 0 0 0 1 0
box 0 0 29072 45152
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
