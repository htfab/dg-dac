magic
tech sky130A
magscale 1 2
timestamp 1748333645
<< pwell >>
rect -2911 -1511 2911 1511
<< mvpsubdiff >>
rect -2845 1433 2845 1445
rect -2845 1399 -2737 1433
rect 2737 1399 2845 1433
rect -2845 1387 2845 1399
rect -2845 1337 -2787 1387
rect -2845 -1337 -2833 1337
rect -2799 -1337 -2787 1337
rect 2787 1337 2845 1387
rect -2845 -1387 -2787 -1337
rect 2787 -1337 2799 1337
rect 2833 -1337 2845 1337
rect 2787 -1387 2845 -1337
rect -2845 -1399 2845 -1387
rect -2845 -1433 -2737 -1399
rect 2737 -1433 2845 -1399
rect -2845 -1445 2845 -1433
<< mvpsubdiffcont >>
rect -2737 1399 2737 1433
rect -2833 -1337 -2799 1337
rect 2799 -1337 2833 1337
rect -2737 -1433 2737 -1399
<< xpolycontact >>
rect -2691 859 -2621 1291
rect -2691 -1291 -2621 -859
rect -2525 859 -2455 1291
rect -2525 -1291 -2455 -859
rect -2359 859 -2289 1291
rect -2359 -1291 -2289 -859
rect -2193 859 -2123 1291
rect -2193 -1291 -2123 -859
rect -2027 859 -1957 1291
rect -2027 -1291 -1957 -859
rect -1861 859 -1791 1291
rect -1861 -1291 -1791 -859
rect -1695 859 -1625 1291
rect -1695 -1291 -1625 -859
rect -1529 859 -1459 1291
rect -1529 -1291 -1459 -859
rect -1363 859 -1293 1291
rect -1363 -1291 -1293 -859
rect -1197 859 -1127 1291
rect -1197 -1291 -1127 -859
rect -1031 859 -961 1291
rect -1031 -1291 -961 -859
rect -865 859 -795 1291
rect -865 -1291 -795 -859
rect -699 859 -629 1291
rect -699 -1291 -629 -859
rect -533 859 -463 1291
rect -533 -1291 -463 -859
rect -367 859 -297 1291
rect -367 -1291 -297 -859
rect -201 859 -131 1291
rect -201 -1291 -131 -859
rect -35 859 35 1291
rect -35 -1291 35 -859
rect 131 859 201 1291
rect 131 -1291 201 -859
rect 297 859 367 1291
rect 297 -1291 367 -859
rect 463 859 533 1291
rect 463 -1291 533 -859
rect 629 859 699 1291
rect 629 -1291 699 -859
rect 795 859 865 1291
rect 795 -1291 865 -859
rect 961 859 1031 1291
rect 961 -1291 1031 -859
rect 1127 859 1197 1291
rect 1127 -1291 1197 -859
rect 1293 859 1363 1291
rect 1293 -1291 1363 -859
rect 1459 859 1529 1291
rect 1459 -1291 1529 -859
rect 1625 859 1695 1291
rect 1625 -1291 1695 -859
rect 1791 859 1861 1291
rect 1791 -1291 1861 -859
rect 1957 859 2027 1291
rect 1957 -1291 2027 -859
rect 2123 859 2193 1291
rect 2123 -1291 2193 -859
rect 2289 859 2359 1291
rect 2289 -1291 2359 -859
rect 2455 859 2525 1291
rect 2455 -1291 2525 -859
rect 2621 859 2691 1291
rect 2621 -1291 2691 -859
<< xpolyres >>
rect -2691 -859 -2621 859
rect -2525 -859 -2455 859
rect -2359 -859 -2289 859
rect -2193 -859 -2123 859
rect -2027 -859 -1957 859
rect -1861 -859 -1791 859
rect -1695 -859 -1625 859
rect -1529 -859 -1459 859
rect -1363 -859 -1293 859
rect -1197 -859 -1127 859
rect -1031 -859 -961 859
rect -865 -859 -795 859
rect -699 -859 -629 859
rect -533 -859 -463 859
rect -367 -859 -297 859
rect -201 -859 -131 859
rect -35 -859 35 859
rect 131 -859 201 859
rect 297 -859 367 859
rect 463 -859 533 859
rect 629 -859 699 859
rect 795 -859 865 859
rect 961 -859 1031 859
rect 1127 -859 1197 859
rect 1293 -859 1363 859
rect 1459 -859 1529 859
rect 1625 -859 1695 859
rect 1791 -859 1861 859
rect 1957 -859 2027 859
rect 2123 -859 2193 859
rect 2289 -859 2359 859
rect 2455 -859 2525 859
rect 2621 -859 2691 859
<< locali >>
rect -2833 1399 -2737 1433
rect 2737 1399 2833 1433
rect -2833 1337 -2799 1399
rect 2799 1337 2833 1399
rect -2833 -1399 -2799 -1337
rect 2799 -1399 2833 -1337
rect -2833 -1433 -2737 -1399
rect 2737 -1433 2833 -1399
<< viali >>
rect -2675 876 -2637 1273
rect -2509 876 -2471 1273
rect -2343 876 -2305 1273
rect -2177 876 -2139 1273
rect -2011 876 -1973 1273
rect -1845 876 -1807 1273
rect -1679 876 -1641 1273
rect -1513 876 -1475 1273
rect -1347 876 -1309 1273
rect -1181 876 -1143 1273
rect -1015 876 -977 1273
rect -849 876 -811 1273
rect -683 876 -645 1273
rect -517 876 -479 1273
rect -351 876 -313 1273
rect -185 876 -147 1273
rect -19 876 19 1273
rect 147 876 185 1273
rect 313 876 351 1273
rect 479 876 517 1273
rect 645 876 683 1273
rect 811 876 849 1273
rect 977 876 1015 1273
rect 1143 876 1181 1273
rect 1309 876 1347 1273
rect 1475 876 1513 1273
rect 1641 876 1679 1273
rect 1807 876 1845 1273
rect 1973 876 2011 1273
rect 2139 876 2177 1273
rect 2305 876 2343 1273
rect 2471 876 2509 1273
rect 2637 876 2675 1273
rect -2675 -1273 -2637 -876
rect -2509 -1273 -2471 -876
rect -2343 -1273 -2305 -876
rect -2177 -1273 -2139 -876
rect -2011 -1273 -1973 -876
rect -1845 -1273 -1807 -876
rect -1679 -1273 -1641 -876
rect -1513 -1273 -1475 -876
rect -1347 -1273 -1309 -876
rect -1181 -1273 -1143 -876
rect -1015 -1273 -977 -876
rect -849 -1273 -811 -876
rect -683 -1273 -645 -876
rect -517 -1273 -479 -876
rect -351 -1273 -313 -876
rect -185 -1273 -147 -876
rect -19 -1273 19 -876
rect 147 -1273 185 -876
rect 313 -1273 351 -876
rect 479 -1273 517 -876
rect 645 -1273 683 -876
rect 811 -1273 849 -876
rect 977 -1273 1015 -876
rect 1143 -1273 1181 -876
rect 1309 -1273 1347 -876
rect 1475 -1273 1513 -876
rect 1641 -1273 1679 -876
rect 1807 -1273 1845 -876
rect 1973 -1273 2011 -876
rect 2139 -1273 2177 -876
rect 2305 -1273 2343 -876
rect 2471 -1273 2509 -876
rect 2637 -1273 2675 -876
<< metal1 >>
rect -2681 1273 -2631 1285
rect -2681 876 -2675 1273
rect -2637 876 -2631 1273
rect -2681 864 -2631 876
rect -2515 1273 -2465 1285
rect -2515 876 -2509 1273
rect -2471 876 -2465 1273
rect -2515 864 -2465 876
rect -2349 1273 -2299 1285
rect -2349 876 -2343 1273
rect -2305 876 -2299 1273
rect -2349 864 -2299 876
rect -2183 1273 -2133 1285
rect -2183 876 -2177 1273
rect -2139 876 -2133 1273
rect -2183 864 -2133 876
rect -2017 1273 -1967 1285
rect -2017 876 -2011 1273
rect -1973 876 -1967 1273
rect -2017 864 -1967 876
rect -1851 1273 -1801 1285
rect -1851 876 -1845 1273
rect -1807 876 -1801 1273
rect -1851 864 -1801 876
rect -1685 1273 -1635 1285
rect -1685 876 -1679 1273
rect -1641 876 -1635 1273
rect -1685 864 -1635 876
rect -1519 1273 -1469 1285
rect -1519 876 -1513 1273
rect -1475 876 -1469 1273
rect -1519 864 -1469 876
rect -1353 1273 -1303 1285
rect -1353 876 -1347 1273
rect -1309 876 -1303 1273
rect -1353 864 -1303 876
rect -1187 1273 -1137 1285
rect -1187 876 -1181 1273
rect -1143 876 -1137 1273
rect -1187 864 -1137 876
rect -1021 1273 -971 1285
rect -1021 876 -1015 1273
rect -977 876 -971 1273
rect -1021 864 -971 876
rect -855 1273 -805 1285
rect -855 876 -849 1273
rect -811 876 -805 1273
rect -855 864 -805 876
rect -689 1273 -639 1285
rect -689 876 -683 1273
rect -645 876 -639 1273
rect -689 864 -639 876
rect -523 1273 -473 1285
rect -523 876 -517 1273
rect -479 876 -473 1273
rect -523 864 -473 876
rect -357 1273 -307 1285
rect -357 876 -351 1273
rect -313 876 -307 1273
rect -357 864 -307 876
rect -191 1273 -141 1285
rect -191 876 -185 1273
rect -147 876 -141 1273
rect -191 864 -141 876
rect -25 1273 25 1285
rect -25 876 -19 1273
rect 19 876 25 1273
rect -25 864 25 876
rect 141 1273 191 1285
rect 141 876 147 1273
rect 185 876 191 1273
rect 141 864 191 876
rect 307 1273 357 1285
rect 307 876 313 1273
rect 351 876 357 1273
rect 307 864 357 876
rect 473 1273 523 1285
rect 473 876 479 1273
rect 517 876 523 1273
rect 473 864 523 876
rect 639 1273 689 1285
rect 639 876 645 1273
rect 683 876 689 1273
rect 639 864 689 876
rect 805 1273 855 1285
rect 805 876 811 1273
rect 849 876 855 1273
rect 805 864 855 876
rect 971 1273 1021 1285
rect 971 876 977 1273
rect 1015 876 1021 1273
rect 971 864 1021 876
rect 1137 1273 1187 1285
rect 1137 876 1143 1273
rect 1181 876 1187 1273
rect 1137 864 1187 876
rect 1303 1273 1353 1285
rect 1303 876 1309 1273
rect 1347 876 1353 1273
rect 1303 864 1353 876
rect 1469 1273 1519 1285
rect 1469 876 1475 1273
rect 1513 876 1519 1273
rect 1469 864 1519 876
rect 1635 1273 1685 1285
rect 1635 876 1641 1273
rect 1679 876 1685 1273
rect 1635 864 1685 876
rect 1801 1273 1851 1285
rect 1801 876 1807 1273
rect 1845 876 1851 1273
rect 1801 864 1851 876
rect 1967 1273 2017 1285
rect 1967 876 1973 1273
rect 2011 876 2017 1273
rect 1967 864 2017 876
rect 2133 1273 2183 1285
rect 2133 876 2139 1273
rect 2177 876 2183 1273
rect 2133 864 2183 876
rect 2299 1273 2349 1285
rect 2299 876 2305 1273
rect 2343 876 2349 1273
rect 2299 864 2349 876
rect 2465 1273 2515 1285
rect 2465 876 2471 1273
rect 2509 876 2515 1273
rect 2465 864 2515 876
rect 2631 1273 2681 1285
rect 2631 876 2637 1273
rect 2675 876 2681 1273
rect 2631 864 2681 876
rect -2681 -876 -2631 -864
rect -2681 -1273 -2675 -876
rect -2637 -1273 -2631 -876
rect -2681 -1285 -2631 -1273
rect -2515 -876 -2465 -864
rect -2515 -1273 -2509 -876
rect -2471 -1273 -2465 -876
rect -2515 -1285 -2465 -1273
rect -2349 -876 -2299 -864
rect -2349 -1273 -2343 -876
rect -2305 -1273 -2299 -876
rect -2349 -1285 -2299 -1273
rect -2183 -876 -2133 -864
rect -2183 -1273 -2177 -876
rect -2139 -1273 -2133 -876
rect -2183 -1285 -2133 -1273
rect -2017 -876 -1967 -864
rect -2017 -1273 -2011 -876
rect -1973 -1273 -1967 -876
rect -2017 -1285 -1967 -1273
rect -1851 -876 -1801 -864
rect -1851 -1273 -1845 -876
rect -1807 -1273 -1801 -876
rect -1851 -1285 -1801 -1273
rect -1685 -876 -1635 -864
rect -1685 -1273 -1679 -876
rect -1641 -1273 -1635 -876
rect -1685 -1285 -1635 -1273
rect -1519 -876 -1469 -864
rect -1519 -1273 -1513 -876
rect -1475 -1273 -1469 -876
rect -1519 -1285 -1469 -1273
rect -1353 -876 -1303 -864
rect -1353 -1273 -1347 -876
rect -1309 -1273 -1303 -876
rect -1353 -1285 -1303 -1273
rect -1187 -876 -1137 -864
rect -1187 -1273 -1181 -876
rect -1143 -1273 -1137 -876
rect -1187 -1285 -1137 -1273
rect -1021 -876 -971 -864
rect -1021 -1273 -1015 -876
rect -977 -1273 -971 -876
rect -1021 -1285 -971 -1273
rect -855 -876 -805 -864
rect -855 -1273 -849 -876
rect -811 -1273 -805 -876
rect -855 -1285 -805 -1273
rect -689 -876 -639 -864
rect -689 -1273 -683 -876
rect -645 -1273 -639 -876
rect -689 -1285 -639 -1273
rect -523 -876 -473 -864
rect -523 -1273 -517 -876
rect -479 -1273 -473 -876
rect -523 -1285 -473 -1273
rect -357 -876 -307 -864
rect -357 -1273 -351 -876
rect -313 -1273 -307 -876
rect -357 -1285 -307 -1273
rect -191 -876 -141 -864
rect -191 -1273 -185 -876
rect -147 -1273 -141 -876
rect -191 -1285 -141 -1273
rect -25 -876 25 -864
rect -25 -1273 -19 -876
rect 19 -1273 25 -876
rect -25 -1285 25 -1273
rect 141 -876 191 -864
rect 141 -1273 147 -876
rect 185 -1273 191 -876
rect 141 -1285 191 -1273
rect 307 -876 357 -864
rect 307 -1273 313 -876
rect 351 -1273 357 -876
rect 307 -1285 357 -1273
rect 473 -876 523 -864
rect 473 -1273 479 -876
rect 517 -1273 523 -876
rect 473 -1285 523 -1273
rect 639 -876 689 -864
rect 639 -1273 645 -876
rect 683 -1273 689 -876
rect 639 -1285 689 -1273
rect 805 -876 855 -864
rect 805 -1273 811 -876
rect 849 -1273 855 -876
rect 805 -1285 855 -1273
rect 971 -876 1021 -864
rect 971 -1273 977 -876
rect 1015 -1273 1021 -876
rect 971 -1285 1021 -1273
rect 1137 -876 1187 -864
rect 1137 -1273 1143 -876
rect 1181 -1273 1187 -876
rect 1137 -1285 1187 -1273
rect 1303 -876 1353 -864
rect 1303 -1273 1309 -876
rect 1347 -1273 1353 -876
rect 1303 -1285 1353 -1273
rect 1469 -876 1519 -864
rect 1469 -1273 1475 -876
rect 1513 -1273 1519 -876
rect 1469 -1285 1519 -1273
rect 1635 -876 1685 -864
rect 1635 -1273 1641 -876
rect 1679 -1273 1685 -876
rect 1635 -1285 1685 -1273
rect 1801 -876 1851 -864
rect 1801 -1273 1807 -876
rect 1845 -1273 1851 -876
rect 1801 -1285 1851 -1273
rect 1967 -876 2017 -864
rect 1967 -1273 1973 -876
rect 2011 -1273 2017 -876
rect 1967 -1285 2017 -1273
rect 2133 -876 2183 -864
rect 2133 -1273 2139 -876
rect 2177 -1273 2183 -876
rect 2133 -1285 2183 -1273
rect 2299 -876 2349 -864
rect 2299 -1273 2305 -876
rect 2343 -1273 2349 -876
rect 2299 -1285 2349 -1273
rect 2465 -876 2515 -864
rect 2465 -1273 2471 -876
rect 2509 -1273 2515 -876
rect 2465 -1285 2515 -1273
rect 2631 -876 2681 -864
rect 2631 -1273 2637 -876
rect 2675 -1273 2681 -876
rect 2631 -1285 2681 -1273
<< properties >>
string FIXED_BBOX -2816 -1416 2816 1416
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 8.75 m 1 nx 33 wmin 0.350 lmin 0.50 class resistor rho 2000 val 51.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
