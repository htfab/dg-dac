magic
tech sky130A
magscale 1 2
timestamp 1748338180
<< dnwell >>
rect 5459 12246 22267 32915
<< nwell >>
rect 5349 32709 22377 33025
rect 5349 12452 5665 32709
rect 22061 12452 22377 32709
rect 5349 12136 22377 12452
<< mvnsubdiff >>
rect 5416 32938 22310 32958
rect 5416 32904 5496 32938
rect 22230 32904 22310 32938
rect 5416 32884 22310 32904
rect 5416 32878 5490 32884
rect 5416 12283 5436 32878
rect 5470 12283 5490 32878
rect 5416 12277 5490 12283
rect 22236 32878 22310 32884
rect 22236 12283 22256 32878
rect 22290 12283 22310 32878
rect 22236 12277 22310 12283
rect 5416 12257 22310 12277
rect 5416 12223 5496 12257
rect 22230 12223 22310 12257
rect 5416 12203 22310 12223
<< mvnsubdiffcont >>
rect 5496 32904 22230 32938
rect 5436 12283 5470 32878
rect 22256 12283 22290 32878
rect 5496 12223 22230 12257
<< locali >>
rect 5436 32904 5496 32938
rect 22230 32904 22290 32938
rect 5436 32878 5470 32904
rect 5436 12257 5470 12283
rect 22256 32878 22290 32904
rect 22256 12257 22290 12283
rect 5436 12223 5496 12257
rect 22230 12223 22290 12257
use toplevel  toplevel_0
timestamp 1748338119
transform 1 0 0 0 1 0
box 0 0 29072 45152
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
