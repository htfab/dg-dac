magic
tech sky130A
magscale 1 2
timestamp 1748318706
<< metal1 >>
rect -264 4657 -204 4663
rect 13544 4657 13604 4663
rect -204 4598 13544 4656
rect -264 4591 -204 4597
rect 13544 4591 13604 4597
rect 3694 3562 3728 4551
rect 6390 3562 6424 4551
rect 9086 3562 9120 4551
rect 9591 3908 9625 4113
rect 11482 3556 11516 4557
rect 11782 3562 11816 4551
rect -564 3525 -504 3531
rect 13844 3525 13904 3531
rect -504 3466 13844 3524
rect -564 3459 -504 3465
rect 13844 3459 13904 3465
rect 8177 3387 8229 3393
rect 2785 3381 2837 3387
rect 4442 3381 4494 3387
rect 2837 3335 4442 3369
rect 2785 3323 2837 3329
rect 4494 3335 8177 3369
rect 10873 3378 10925 3384
rect 8229 3335 10873 3369
rect 8177 3329 8229 3335
rect 4442 3323 4494 3329
rect 10873 3320 10925 3326
<< via1 >>
rect -264 4597 -204 4657
rect 13544 4597 13604 4657
rect -564 3465 -504 3525
rect 13844 3465 13904 3525
rect 2785 3329 2837 3381
rect 4442 3329 4494 3381
rect 8177 3335 8229 3387
rect 10873 3326 10925 3378
<< metal2 >>
rect -270 4597 -264 4657
rect -204 4597 -198 4657
rect 13538 4597 13544 4657
rect 13604 4597 13610 4657
rect -570 3465 -564 3525
rect -504 3465 -498 3525
rect -564 2785 -504 3465
rect -571 2729 -562 2785
rect -506 2729 -497 2785
rect -564 2185 -504 2729
rect -264 2485 -204 4597
rect 1503 3301 1537 4113
rect 2794 3381 2828 4021
rect 2779 3329 2785 3381
rect 2837 3329 2843 3381
rect 4199 3369 4233 4113
rect 5490 3446 5524 4021
rect 4451 3412 5524 3446
rect 4451 3381 4485 3412
rect 3186 3335 4233 3369
rect 3186 3301 3220 3335
rect 4436 3329 4442 3381
rect 4494 3329 4500 3381
rect 6895 3369 6929 4113
rect 8186 3387 8220 4021
rect 4528 3335 6929 3369
rect 8171 3335 8177 3387
rect 8229 3335 8235 3387
rect 4528 3301 4562 3335
rect 9591 3301 9625 4095
rect 10882 3378 10916 4021
rect 10867 3326 10873 3378
rect 10925 3326 10931 3378
rect 579 3267 1537 3301
rect 1921 3267 3220 3301
rect 3263 3267 4562 3301
rect 4605 3267 9625 3301
rect 207 2787 263 2794
rect 205 2785 265 2787
rect 205 2729 207 2785
rect 263 2729 265 2785
rect 205 2672 265 2729
rect 13544 2485 13604 4597
rect 13838 3465 13844 3525
rect 13904 3465 13910 3525
rect 13844 2785 13904 3465
rect 13837 2729 13846 2785
rect 13902 2729 13911 2785
rect -271 2429 -262 2485
rect -206 2429 -197 2485
rect 13537 2429 13546 2485
rect 13602 2429 13611 2485
rect -571 2129 -562 2185
rect -506 2129 -497 2185
rect -564 1585 -504 2129
rect -264 1885 -204 2429
rect 13544 1885 13604 2429
rect 13844 2185 13904 2729
rect 13837 2129 13846 2185
rect 13902 2129 13911 2185
rect -271 1829 -262 1885
rect -206 1829 -197 1885
rect 13537 1829 13546 1885
rect 13602 1829 13611 1885
rect -571 1529 -562 1585
rect -506 1529 -497 1585
rect -564 985 -504 1529
rect -264 1285 -204 1829
rect 13544 1285 13604 1829
rect 13844 1585 13904 2129
rect 13837 1529 13846 1585
rect 13902 1529 13911 1585
rect -271 1229 -262 1285
rect -206 1229 -197 1285
rect 13537 1229 13546 1285
rect 13602 1229 13611 1285
rect -571 929 -562 985
rect -506 929 -497 985
rect -564 385 -504 929
rect -264 685 -204 1229
rect 13544 685 13604 1229
rect 13844 985 13904 1529
rect 13837 929 13846 985
rect 13902 929 13911 985
rect -271 629 -262 685
rect -206 629 -197 685
rect 13537 629 13546 685
rect 13602 629 13611 685
rect -264 627 -204 629
rect 13544 627 13604 629
rect 13844 385 13904 929
rect -571 329 -562 385
rect -506 329 -497 385
rect 13837 329 13846 385
rect 13902 329 13911 385
rect -564 327 -504 329
rect 13844 327 13904 329
rect 3263 78 3297 224
rect 3960 78 3994 224
rect 4605 78 4639 224
rect 5302 78 5336 224
rect 5947 78 5981 224
rect 6644 78 6678 224
rect 7289 78 7323 224
rect 7986 78 8020 224
rect 8631 78 8665 224
rect 9328 78 9362 224
rect 9973 78 10007 224
rect 10670 78 10704 224
rect 11315 78 11349 224
rect 12012 78 12046 224
rect 12657 78 12691 224
rect 13354 78 13388 224
<< via2 >>
rect -562 2729 -506 2785
rect 207 2729 263 2785
rect 13846 2729 13902 2785
rect -262 2429 -206 2485
rect 13546 2429 13602 2485
rect -562 2129 -506 2185
rect 13846 2129 13902 2185
rect -262 1829 -206 1885
rect 13546 1829 13602 1885
rect -562 1529 -506 1585
rect 13846 1529 13902 1585
rect -262 1229 -206 1285
rect 13546 1229 13602 1285
rect -562 929 -506 985
rect 13846 929 13902 985
rect -262 629 -206 685
rect 13546 629 13602 685
rect -562 329 -506 385
rect 13846 329 13902 385
<< metal3 >>
rect -567 2787 -501 2790
rect 202 2787 268 2790
rect 13841 2787 13907 2790
rect -567 2785 13907 2787
rect -567 2729 -562 2785
rect -506 2729 207 2785
rect 263 2729 13846 2785
rect 13902 2729 13907 2785
rect -567 2727 13907 2729
rect -567 2724 -501 2727
rect 202 2724 268 2727
rect 13841 2724 13907 2727
rect -267 2487 -201 2490
rect 13541 2487 13607 2490
rect -267 2485 13607 2487
rect -267 2429 -262 2485
rect -206 2429 13546 2485
rect 13602 2429 13607 2485
rect -267 2427 13607 2429
rect -267 2424 -201 2427
rect 13541 2424 13607 2427
rect -567 2187 -501 2190
rect 13841 2187 13907 2190
rect -567 2185 13907 2187
rect -567 2129 -562 2185
rect -506 2129 13846 2185
rect 13902 2129 13907 2185
rect -567 2127 13907 2129
rect -567 2124 -501 2127
rect 13841 2124 13907 2127
rect -267 1887 -201 1890
rect 13541 1887 13607 1890
rect -267 1885 13607 1887
rect -267 1829 -262 1885
rect -206 1829 13546 1885
rect 13602 1829 13607 1885
rect -267 1827 13607 1829
rect -267 1824 -201 1827
rect 13541 1824 13607 1827
rect -567 1587 -501 1590
rect 13841 1587 13907 1590
rect -567 1585 13907 1587
rect -567 1529 -562 1585
rect -506 1529 13846 1585
rect 13902 1529 13907 1585
rect -567 1527 13907 1529
rect -567 1524 -501 1527
rect 13841 1524 13907 1527
rect -267 1287 -201 1290
rect 13541 1287 13607 1290
rect -267 1285 13607 1287
rect -267 1229 -262 1285
rect -206 1229 13546 1285
rect 13602 1229 13607 1285
rect -267 1227 13607 1229
rect -267 1224 -201 1227
rect 13541 1224 13607 1227
rect -567 987 -501 990
rect 13841 987 13907 990
rect -567 985 13907 987
rect -567 929 -562 985
rect -506 929 13846 985
rect 13902 929 13907 985
rect -567 927 13907 929
rect -567 924 -501 927
rect 13841 924 13907 927
rect -267 687 -201 690
rect 13541 687 13607 690
rect -267 685 13607 687
rect -267 629 -262 685
rect -206 629 13546 685
rect 13602 629 13607 685
rect -267 627 13607 629
rect -267 624 -201 627
rect 13541 624 13607 627
rect -567 387 -501 390
rect 13841 387 13907 390
rect -567 385 13907 387
rect -567 329 -562 385
rect -506 329 13846 385
rect 13902 329 13907 385
rect -567 327 13907 329
rect -567 324 -501 327
rect 13841 324 13907 327
use decoder4  decoder4_0
timestamp 1748318706
transform 0 1 0 -1 0 2996
box -305 0 2996 13410
use xor2  xor2_0
array 0 3 2696 0 0 1292
timestamp 1748318706
transform -1 0 12097 0 -1 4692
box 0 0 2696 1292
<< labels >>
flabel metal2 3960 78 3994 224 0 FreeSans 128 90 0 0 D[0]
port 10 nsew signal output
flabel metal2 3263 78 3297 224 0 FreeSans 128 90 0 0 D[1]
port 6 nsew signal output
flabel metal2 5302 78 5336 224 0 FreeSans 128 90 0 0 D[2]
port 4 nsew signal output
flabel metal2 4605 78 4639 224 0 FreeSans 128 90 0 0 D[3]
port 2 nsew signal output
flabel metal2 6644 78 6678 224 0 FreeSans 128 90 0 0 D[4]
port 20 nsew signal output
flabel metal2 5947 78 5981 224 0 FreeSans 128 90 0 0 D[5]
port 18 nsew signal output
flabel metal2 7986 78 8020 224 0 FreeSans 128 90 0 0 D[6]
port 16 nsew signal output
flabel metal2 7289 78 7323 224 0 FreeSans 128 90 0 0 D[7]
port 14 nsew signal output
flabel metal2 9328 78 9362 224 0 FreeSans 128 90 0 0 D[8]
port 8 nsew signal output
flabel metal2 8631 78 8665 224 0 FreeSans 128 90 0 0 D[9]
port 5 nsew signal output
flabel metal2 10670 78 10704 224 0 FreeSans 128 90 0 0 D[10]
port 3 nsew signal output
flabel metal2 9973 78 10007 224 0 FreeSans 128 90 0 0 D[11]
port 1 nsew signal output
flabel metal2 12012 78 12046 224 0 FreeSans 128 90 0 0 D[12]
port 19 nsew signal output
flabel metal2 11315 78 11349 224 0 FreeSans 128 90 0 0 D[13]
port 17 nsew signal output
flabel metal2 13354 78 13388 224 0 FreeSans 128 90 0 0 D[14]
port 15 nsew signal output
flabel metal2 12657 78 12691 224 0 FreeSans 128 90 0 0 D[15]
port 12 nsew signal output
flabel metal3 36 2727 13304 2787 0 FreeSans 128 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal3 36 2427 13304 2487 0 FreeSans 128 90 0 0 VSS
port 21 nsew ground bidirectional
flabel metal1 9086 3562 9120 4551 0 FreeSans 256 0 0 0 IN[0]
port 22 nsew signal input
flabel metal1 11782 3562 11816 4551 0 FreeSans 256 0 0 0 IN[1]
port 23 nsew signal input
flabel metal1 3694 3562 3728 4551 0 FreeSans 256 0 0 0 IN[2]
port 24 nsew signal input
flabel metal1 6390 3562 6424 4551 0 FreeSans 256 0 0 0 IN[3]
port 25 nsew signal input
flabel metal1 11482 3556 11516 4557 0 FreeSans 256 0 0 0 IN[4]
port 26 nsew signal input
<< end >>
