magic
tech sky130A
magscale 1 2
timestamp 1740620545
<< locali >>
rect 150 7058 250 7070
rect 150 6466 156 7058
rect 244 6466 250 7058
rect 150 6454 250 6466
rect 5572 7058 5672 7070
rect 5572 6466 5578 7058
rect 5666 6466 5672 7058
rect 5572 6454 5672 6466
rect 150 6074 253 6086
rect 150 5324 156 6074
rect 244 5324 253 6074
rect 150 5312 253 5324
rect 5572 6074 5672 6086
rect 5572 5324 5578 6074
rect 5666 5324 5672 6074
rect 5572 5312 5672 5324
rect 0 4932 112 4944
rect 0 2282 6 4932
rect 106 2282 112 4932
rect 0 2270 112 2282
rect 5710 4932 5822 4944
rect 5710 2282 5716 4932
rect 5816 2282 5822 4932
rect 5710 2270 5822 2282
rect 150 1890 253 1902
rect 150 1140 156 1890
rect 244 1140 253 1890
rect 150 1128 253 1140
rect 5572 1890 5672 1902
rect 5572 1140 5578 1890
rect 5666 1140 5672 1890
rect 5572 1128 5672 1140
rect 150 748 250 760
rect 150 156 156 748
rect 244 156 250 748
rect 150 144 250 156
rect 5572 748 5672 760
rect 5572 156 5578 748
rect 5666 156 5672 748
rect 5572 144 5672 156
<< viali >>
rect 156 6466 244 7058
rect 5578 6466 5666 7058
rect 156 5324 244 6074
rect 5578 5324 5666 6074
rect 6 2282 106 4932
rect 5716 2282 5816 4932
rect 156 1140 244 1890
rect 5578 1140 5666 1890
rect 156 156 244 748
rect 5578 156 5666 748
<< metal1 >>
rect 0 7058 250 7070
rect 0 6466 6 7058
rect 94 6466 156 7058
rect 244 6466 250 7058
rect 0 6454 250 6466
rect 5572 7058 5822 7070
rect 5572 6466 5578 7058
rect 5666 6466 5728 7058
rect 5816 6466 5822 7058
rect 5572 6454 5822 6466
rect 150 6074 250 6086
rect 150 5324 156 6074
rect 244 5324 250 6074
rect 150 5312 250 5324
rect 5572 6074 5672 6086
rect 5572 5324 5578 6074
rect 5666 5324 5672 6074
rect 5572 5312 5672 5324
rect 0 4932 112 4944
rect 0 2282 6 4932
rect 106 4898 112 4932
rect 5710 4932 5822 4944
rect 5710 4898 5716 4932
rect 106 4717 456 4898
rect 106 4647 386 4717
rect 106 4466 456 4647
rect 552 4717 788 4898
rect 552 4647 635 4717
rect 705 4647 788 4717
rect 552 4466 788 4647
rect 884 4717 1120 4898
rect 884 4647 967 4717
rect 1037 4647 1120 4717
rect 884 4466 1120 4647
rect 1216 4717 1452 4898
rect 1216 4647 1299 4717
rect 1369 4647 1452 4717
rect 1216 4466 1452 4647
rect 1548 4717 1784 4898
rect 1548 4647 1631 4717
rect 1701 4647 1784 4717
rect 1548 4466 1784 4647
rect 1880 4717 2116 4898
rect 1880 4647 1963 4717
rect 2033 4647 2116 4717
rect 1880 4466 2116 4647
rect 2212 4717 2448 4898
rect 2212 4647 2295 4717
rect 2365 4647 2448 4717
rect 2212 4466 2448 4647
rect 2544 4717 2780 4898
rect 2544 4647 2627 4717
rect 2697 4647 2780 4717
rect 2544 4466 2780 4647
rect 106 2748 112 4466
rect 2876 3382 2946 4898
rect 3042 4422 3112 4898
rect 3208 4717 3444 4898
rect 3208 4647 3291 4717
rect 3361 4647 3444 4717
rect 3208 4466 3444 4647
rect 3540 4717 3776 4898
rect 3540 4647 3623 4717
rect 3693 4647 3776 4717
rect 3540 4466 3776 4647
rect 3872 4717 4108 4898
rect 3872 4647 3955 4717
rect 4025 4647 4108 4717
rect 3872 4466 4108 4647
rect 4204 4717 4440 4898
rect 4204 4647 4287 4717
rect 4357 4647 4440 4717
rect 4204 4466 4440 4647
rect 4536 4717 4772 4898
rect 4536 4647 4619 4717
rect 4689 4647 4772 4717
rect 4536 4466 4772 4647
rect 4868 4717 5104 4898
rect 4868 4647 4951 4717
rect 5021 4647 5104 4717
rect 4868 4466 5104 4647
rect 5200 4717 5436 4898
rect 5200 4647 5283 4717
rect 5353 4647 5436 4717
rect 5200 4466 5436 4647
rect 5532 4466 5716 4898
rect 3042 4346 3112 4352
rect 2870 3312 2876 3382
rect 2946 3312 2952 3382
rect 5710 2748 5716 4466
rect 106 2316 290 2748
rect 386 2567 622 2748
rect 386 2497 469 2567
rect 539 2497 622 2567
rect 386 2316 622 2497
rect 718 2567 954 2748
rect 718 2497 801 2567
rect 871 2497 954 2567
rect 718 2316 954 2497
rect 1050 2567 1286 2748
rect 1050 2497 1133 2567
rect 1203 2497 1286 2567
rect 1050 2316 1286 2497
rect 1382 2567 1618 2748
rect 1382 2497 1465 2567
rect 1535 2497 1618 2567
rect 1382 2316 1618 2497
rect 1714 2567 1950 2748
rect 1714 2497 1797 2567
rect 1867 2497 1950 2567
rect 1714 2316 1950 2497
rect 2046 2567 2282 2748
rect 2046 2497 2129 2567
rect 2199 2497 2282 2567
rect 2046 2316 2282 2497
rect 2378 2567 2614 2748
rect 2378 2497 2461 2567
rect 2531 2497 2614 2567
rect 2378 2316 2614 2497
rect 2710 2567 2946 2748
rect 2710 2497 2793 2567
rect 2863 2497 2946 2567
rect 2710 2316 2946 2497
rect 3042 2567 3278 2748
rect 3042 2497 3125 2567
rect 3195 2497 3278 2567
rect 3042 2316 3278 2497
rect 3374 2567 3610 2748
rect 3374 2497 3457 2567
rect 3527 2497 3610 2567
rect 3374 2316 3610 2497
rect 3706 2567 3942 2748
rect 3706 2497 3789 2567
rect 3859 2497 3942 2567
rect 3706 2316 3942 2497
rect 4038 2567 4274 2748
rect 4038 2497 4121 2567
rect 4191 2497 4274 2567
rect 4038 2316 4274 2497
rect 4370 2567 4606 2748
rect 4370 2497 4453 2567
rect 4523 2497 4606 2567
rect 4370 2316 4606 2497
rect 4702 2567 4938 2748
rect 4702 2497 4785 2567
rect 4855 2497 4938 2567
rect 4702 2316 4938 2497
rect 5034 2567 5270 2748
rect 5034 2497 5117 2567
rect 5187 2497 5270 2567
rect 5034 2316 5270 2497
rect 5366 2567 5436 2748
rect 5366 2316 5436 2497
rect 5532 2316 5716 2748
rect 106 2282 112 2316
rect 0 2270 112 2282
rect 5710 2282 5716 2316
rect 5816 2282 5822 4932
rect 5710 2270 5822 2282
rect 150 1890 250 1902
rect 150 1140 156 1890
rect 244 1140 250 1890
rect 150 1128 250 1140
rect 5572 1890 5672 1902
rect 5572 1140 5578 1890
rect 5666 1140 5672 1890
rect 5572 1128 5672 1140
rect 0 748 250 760
rect 0 156 6 748
rect 94 156 156 748
rect 244 156 250 748
rect 0 144 250 156
rect 5572 748 5822 760
rect 5572 156 5578 748
rect 5666 156 5728 748
rect 5816 156 5822 748
rect 5572 144 5822 156
<< via1 >>
rect 6 6466 94 7058
rect 5728 6466 5816 7058
rect 156 5324 244 6074
rect 5578 5324 5666 6074
rect 6 2282 94 4932
rect 386 4647 456 4717
rect 635 4647 705 4717
rect 967 4647 1037 4717
rect 1299 4647 1369 4717
rect 1631 4647 1701 4717
rect 1963 4647 2033 4717
rect 2295 4647 2365 4717
rect 2627 4647 2697 4717
rect 3291 4647 3361 4717
rect 3623 4647 3693 4717
rect 3955 4647 4025 4717
rect 4287 4647 4357 4717
rect 4619 4647 4689 4717
rect 4951 4647 5021 4717
rect 5283 4647 5353 4717
rect 3042 4352 3112 4422
rect 2876 3312 2946 3382
rect 469 2497 539 2567
rect 801 2497 871 2567
rect 1133 2497 1203 2567
rect 1465 2497 1535 2567
rect 1797 2497 1867 2567
rect 2129 2497 2199 2567
rect 2461 2497 2531 2567
rect 2793 2497 2863 2567
rect 3125 2497 3195 2567
rect 3457 2497 3527 2567
rect 3789 2497 3859 2567
rect 4121 2497 4191 2567
rect 4453 2497 4523 2567
rect 4785 2497 4855 2567
rect 5117 2497 5187 2567
rect 5366 2497 5436 2567
rect 5728 2282 5816 4932
rect 156 1140 244 1890
rect 5578 1140 5666 1890
rect 6 156 94 748
rect 5728 156 5816 748
<< metal2 >>
rect 0 7058 100 7214
rect 0 6466 6 7058
rect 94 6466 100 7058
rect 0 4932 100 6466
rect 0 2282 6 4932
rect 94 2282 100 4932
rect 0 748 100 2282
rect 0 156 6 748
rect 94 156 100 748
rect 0 0 100 156
rect 150 6074 250 7214
rect 685 6529 823 7172
rect 961 6701 1099 6839
rect 1237 6701 1375 6839
rect 1513 6701 1651 6839
rect 1789 6701 1927 6839
rect 2065 6701 2203 6839
rect 2341 6701 2479 6839
rect 2617 6701 2755 6839
rect 2893 6701 3031 6839
rect 3169 6701 3307 6839
rect 3445 6701 3583 6839
rect 3721 6701 3859 6839
rect 3997 6701 4135 6839
rect 4273 6701 4411 6839
rect 4549 6701 4687 6839
rect 4825 6701 4963 6839
rect 5101 6701 5239 6839
rect 961 6657 1099 6667
rect 961 6539 971 6657
rect 1089 6539 1099 6657
rect 961 6529 1099 6539
rect 1237 6657 1375 6667
rect 1237 6539 1247 6657
rect 1365 6539 1375 6657
rect 1237 6529 1375 6539
rect 1513 6657 1651 6667
rect 1513 6539 1523 6657
rect 1641 6539 1651 6657
rect 1513 6529 1651 6539
rect 1789 6657 1927 6667
rect 1789 6539 1799 6657
rect 1917 6539 1927 6657
rect 1789 6529 1927 6539
rect 2065 6657 2203 6667
rect 2065 6539 2075 6657
rect 2193 6539 2203 6657
rect 2065 6529 2203 6539
rect 2341 6657 2479 6667
rect 2341 6539 2351 6657
rect 2469 6539 2479 6657
rect 2341 6529 2479 6539
rect 2617 6657 2755 6667
rect 2617 6539 2627 6657
rect 2745 6539 2755 6657
rect 2617 6529 2755 6539
rect 2893 6657 3031 6667
rect 2893 6539 2903 6657
rect 3021 6539 3031 6657
rect 2893 6529 3031 6539
rect 3169 6657 3307 6667
rect 3169 6539 3179 6657
rect 3297 6539 3307 6657
rect 3169 6529 3307 6539
rect 3445 6657 3583 6667
rect 3445 6539 3455 6657
rect 3573 6539 3583 6657
rect 3445 6529 3583 6539
rect 3721 6657 3859 6667
rect 3721 6539 3731 6657
rect 3849 6539 3859 6657
rect 3721 6529 3859 6539
rect 3997 6657 4135 6667
rect 3997 6539 4007 6657
rect 4125 6539 4135 6657
rect 3997 6529 4135 6539
rect 4273 6657 4411 6667
rect 4273 6539 4283 6657
rect 4401 6539 4411 6657
rect 4273 6529 4411 6539
rect 4549 6657 4687 6667
rect 4549 6539 4559 6657
rect 4677 6539 4687 6657
rect 4549 6529 4687 6539
rect 4825 6657 4963 6667
rect 4825 6539 4835 6657
rect 4953 6539 4963 6657
rect 4825 6529 4963 6539
rect 5101 6657 5239 6667
rect 5101 6539 5111 6657
rect 5229 6539 5239 6657
rect 5101 6529 5239 6539
rect 150 5324 156 6074
rect 244 5324 250 6074
rect 5572 6074 5672 7214
rect 583 5613 721 6021
rect 893 5987 963 5996
rect 893 5908 963 5917
rect 1169 5987 1239 5996
rect 1169 5908 1239 5917
rect 1445 5987 1515 5996
rect 1445 5908 1515 5917
rect 1721 5987 1791 5996
rect 1721 5908 1791 5917
rect 1997 5987 2067 5996
rect 1997 5908 2067 5917
rect 2273 5987 2343 5996
rect 2273 5908 2343 5917
rect 2549 5987 2619 5996
rect 2549 5908 2619 5917
rect 2825 5987 2895 5996
rect 2825 5908 2895 5917
rect 3101 5987 3171 5996
rect 3101 5908 3171 5917
rect 3377 5987 3447 5996
rect 3377 5908 3447 5917
rect 3653 5987 3723 5996
rect 3653 5908 3723 5917
rect 3929 5987 3999 5996
rect 3929 5908 3999 5917
rect 4205 5987 4275 5996
rect 4205 5908 4275 5917
rect 4481 5987 4551 5996
rect 4481 5908 4551 5917
rect 4757 5987 4827 5996
rect 4757 5908 4827 5917
rect 5033 5987 5103 5996
rect 5033 5908 5103 5917
rect 150 3377 250 5324
rect 5572 5324 5578 6074
rect 5666 5324 5672 6074
rect 4453 5148 4523 5153
rect 4619 5148 4689 5153
rect 4785 5148 4855 5153
rect 4951 5148 5021 5153
rect 5117 5148 5187 5153
rect 5283 5148 5353 5153
rect 4449 5088 4458 5148
rect 4518 5088 4527 5148
rect 4615 5088 4624 5148
rect 4684 5088 4693 5148
rect 4781 5088 4790 5148
rect 4850 5088 4859 5148
rect 4947 5088 4956 5148
rect 5016 5088 5025 5148
rect 5113 5088 5122 5148
rect 5182 5088 5191 5148
rect 5279 5088 5288 5148
rect 5348 5088 5357 5148
rect 4287 5067 4357 5072
rect 4283 5007 4292 5067
rect 4352 5007 4361 5067
rect 4121 4937 4191 4942
rect 4117 4877 4126 4937
rect 4186 4877 4195 4937
rect 3955 4807 4025 4812
rect 3951 4747 3960 4807
rect 4020 4747 4029 4807
rect 3955 4717 4025 4747
rect 150 3317 155 3377
rect 215 3317 250 3377
rect 150 1890 250 3317
rect 303 4647 386 4717
rect 456 4647 462 4717
rect 629 4647 635 4717
rect 705 4647 711 4717
rect 961 4647 967 4717
rect 1037 4647 1043 4717
rect 1293 4647 1299 4717
rect 1369 4647 1375 4717
rect 1625 4647 1631 4717
rect 1701 4647 1707 4717
rect 1957 4647 1963 4717
rect 2033 4647 2039 4717
rect 2289 4647 2295 4717
rect 2365 4647 2371 4717
rect 2621 4647 2627 4717
rect 2697 4647 2703 4717
rect 3285 4647 3291 4717
rect 3361 4647 3367 4717
rect 3617 4647 3623 4717
rect 3693 4647 3699 4717
rect 3789 4677 3859 4682
rect 303 2126 373 4647
rect 463 2497 469 2567
rect 539 2497 545 2567
rect 469 2126 539 2497
rect 635 2126 705 4647
rect 795 2497 801 2567
rect 871 2497 877 2567
rect 801 2126 871 2497
rect 967 2126 1037 4647
rect 1127 2497 1133 2567
rect 1203 2497 1209 2567
rect 1133 2126 1203 2497
rect 1299 2126 1369 4647
rect 1459 2497 1465 2567
rect 1535 2497 1541 2567
rect 1465 2207 1535 2497
rect 1631 2337 1701 4647
rect 1963 2597 2033 4647
rect 2295 2857 2365 4647
rect 2627 3117 2697 4647
rect 2959 4352 3042 4422
rect 3112 4352 3118 4422
rect 2959 4027 3029 4352
rect 3291 4287 3361 4647
rect 3623 4547 3693 4647
rect 3785 4617 3794 4677
rect 3854 4617 3863 4677
rect 3949 4647 3955 4717
rect 4025 4647 4031 4717
rect 3619 4487 3628 4547
rect 3688 4487 3697 4547
rect 3623 4482 3693 4487
rect 3457 4417 3527 4422
rect 3453 4357 3462 4417
rect 3522 4357 3531 4417
rect 3287 4227 3296 4287
rect 3356 4227 3365 4287
rect 3291 4222 3361 4227
rect 3125 4157 3195 4162
rect 3121 4097 3130 4157
rect 3190 4097 3199 4157
rect 2955 3967 2964 4027
rect 3024 3967 3033 4027
rect 2959 3517 3029 3967
rect 2950 3447 2959 3517
rect 3029 3447 3038 3517
rect 2876 3382 2946 3388
rect 2872 3317 2876 3377
rect 2946 3317 2950 3377
rect 2876 3306 2946 3312
rect 2793 3247 2863 3252
rect 2789 3187 2798 3247
rect 2858 3187 2867 3247
rect 2623 3057 2632 3117
rect 2692 3057 2701 3117
rect 2627 3052 2697 3057
rect 2461 2987 2531 2992
rect 2457 2927 2466 2987
rect 2526 2927 2535 2987
rect 2291 2797 2300 2857
rect 2360 2797 2369 2857
rect 2295 2792 2365 2797
rect 2129 2727 2199 2732
rect 2125 2667 2134 2727
rect 2194 2667 2203 2727
rect 1791 2497 1797 2567
rect 1867 2497 1873 2567
rect 1959 2537 1968 2597
rect 2028 2537 2037 2597
rect 2129 2567 2199 2667
rect 2461 2567 2531 2927
rect 2793 2567 2863 3187
rect 3125 2567 3195 4097
rect 3457 2567 3527 4357
rect 3789 2567 3859 4617
rect 4121 2567 4191 4877
rect 4287 4717 4357 5007
rect 4281 4647 4287 4717
rect 4357 4647 4363 4717
rect 4453 2567 4523 5088
rect 4619 4717 4689 5088
rect 4613 4647 4619 4717
rect 4689 4647 4695 4717
rect 4785 2567 4855 5088
rect 4951 4717 5021 5088
rect 4945 4647 4951 4717
rect 5021 4647 5027 4717
rect 5117 2567 5187 5088
rect 5283 4717 5353 5088
rect 5277 4647 5283 4717
rect 5353 4647 5359 4717
rect 5449 2567 5519 2573
rect 1963 2532 2033 2537
rect 2123 2497 2129 2567
rect 2199 2497 2205 2567
rect 2455 2497 2461 2567
rect 2531 2497 2537 2567
rect 2787 2497 2793 2567
rect 2863 2497 2869 2567
rect 3119 2497 3125 2567
rect 3195 2497 3201 2567
rect 3451 2497 3457 2567
rect 3527 2497 3533 2567
rect 3783 2497 3789 2567
rect 3859 2497 3865 2567
rect 4115 2497 4121 2567
rect 4191 2497 4197 2567
rect 4447 2497 4453 2567
rect 4523 2497 4529 2567
rect 4779 2497 4785 2567
rect 4855 2497 4861 2567
rect 5111 2497 5117 2567
rect 5187 2497 5193 2567
rect 5360 2497 5366 2567
rect 5436 2562 5519 2567
rect 5436 2502 5454 2562
rect 5514 2502 5523 2562
rect 5436 2497 5519 2502
rect 1797 2467 1867 2497
rect 5449 2491 5519 2497
rect 1793 2407 1802 2467
rect 1862 2407 1871 2467
rect 1797 2402 1867 2407
rect 1627 2277 1636 2337
rect 1696 2277 1705 2337
rect 1631 2272 1701 2277
rect 1461 2147 1470 2207
rect 1530 2147 1539 2207
rect 1465 2142 1535 2147
rect 299 2066 308 2126
rect 368 2066 377 2126
rect 465 2066 474 2126
rect 534 2066 543 2126
rect 631 2066 640 2126
rect 700 2066 709 2126
rect 797 2066 806 2126
rect 866 2066 875 2126
rect 963 2066 972 2126
rect 1032 2066 1041 2126
rect 1129 2066 1138 2126
rect 1198 2066 1207 2126
rect 1295 2066 1304 2126
rect 1364 2066 1373 2126
rect 303 2061 373 2066
rect 469 2061 539 2066
rect 635 2061 705 2066
rect 801 2061 871 2066
rect 967 2061 1037 2066
rect 1133 2061 1203 2066
rect 1299 2061 1369 2066
rect 150 1140 156 1890
rect 244 1140 250 1890
rect 5572 1890 5672 5324
rect 719 1297 789 1306
rect 719 1218 789 1227
rect 995 1297 1065 1306
rect 995 1218 1065 1227
rect 1271 1297 1341 1306
rect 1271 1218 1341 1227
rect 1547 1297 1617 1306
rect 1547 1218 1617 1227
rect 1823 1297 1893 1306
rect 1823 1218 1893 1227
rect 2099 1297 2169 1306
rect 2099 1218 2169 1227
rect 2375 1297 2445 1306
rect 2375 1218 2445 1227
rect 2651 1297 2721 1306
rect 2651 1218 2721 1227
rect 2927 1297 2997 1306
rect 2927 1218 2997 1227
rect 3203 1297 3273 1306
rect 3203 1218 3273 1227
rect 3479 1297 3549 1306
rect 3479 1218 3549 1227
rect 3755 1297 3825 1306
rect 3755 1218 3825 1227
rect 4031 1297 4101 1306
rect 4031 1218 4101 1227
rect 4307 1297 4377 1306
rect 4307 1218 4377 1227
rect 4583 1297 4653 1306
rect 4583 1218 4653 1227
rect 4859 1297 4929 1306
rect 4859 1218 4929 1227
rect 5135 1297 5205 1306
rect 5135 1218 5205 1227
rect 150 0 250 1140
rect 5572 1140 5578 1890
rect 5666 1140 5672 1890
rect 583 675 721 685
rect 583 557 593 675
rect 711 557 721 675
rect 583 547 721 557
rect 859 675 997 685
rect 859 557 869 675
rect 987 557 997 675
rect 859 547 997 557
rect 1135 675 1273 685
rect 1135 557 1145 675
rect 1263 557 1273 675
rect 1135 547 1273 557
rect 1411 675 1549 685
rect 1411 557 1421 675
rect 1539 557 1549 675
rect 1411 547 1549 557
rect 1687 675 1825 685
rect 1687 557 1697 675
rect 1815 557 1825 675
rect 1687 547 1825 557
rect 1963 675 2101 685
rect 1963 557 1973 675
rect 2091 557 2101 675
rect 1963 547 2101 557
rect 2239 675 2377 685
rect 2239 557 2249 675
rect 2367 557 2377 675
rect 2239 547 2377 557
rect 2515 675 2653 685
rect 2515 557 2525 675
rect 2643 557 2653 675
rect 2515 547 2653 557
rect 2791 675 2929 685
rect 2791 557 2801 675
rect 2919 557 2929 675
rect 2791 547 2929 557
rect 3067 675 3205 685
rect 3067 557 3077 675
rect 3195 557 3205 675
rect 3067 547 3205 557
rect 3343 675 3481 685
rect 3343 557 3353 675
rect 3471 557 3481 675
rect 3343 547 3481 557
rect 3619 675 3757 685
rect 3619 557 3629 675
rect 3747 557 3757 675
rect 3619 547 3757 557
rect 3895 675 4033 685
rect 3895 557 3905 675
rect 4023 557 4033 675
rect 3895 547 4033 557
rect 4171 675 4309 685
rect 4171 557 4181 675
rect 4299 557 4309 675
rect 4171 547 4309 557
rect 4447 675 4585 685
rect 4447 557 4457 675
rect 4575 557 4585 675
rect 4447 547 4585 557
rect 4723 675 4861 685
rect 4723 557 4733 675
rect 4851 557 4861 675
rect 4723 547 4861 557
rect 4999 675 5137 685
rect 4999 557 5009 675
rect 5127 557 5137 675
rect 4999 547 5137 557
rect 583 375 721 513
rect 859 375 997 513
rect 1135 375 1273 513
rect 1411 375 1549 513
rect 1687 375 1825 513
rect 1963 375 2101 513
rect 2239 375 2377 513
rect 2515 375 2653 513
rect 2791 375 2929 513
rect 3067 375 3205 513
rect 3343 375 3481 513
rect 3619 375 3757 513
rect 3895 375 4033 513
rect 4171 375 4309 513
rect 4447 375 4585 513
rect 4723 375 4861 513
rect 4999 375 5137 513
rect 5572 0 5672 1140
rect 5722 7058 5822 7214
rect 5722 6466 5728 7058
rect 5816 6466 5822 7058
rect 5722 4932 5822 6466
rect 5722 2282 5728 4932
rect 5816 2282 5822 4932
rect 5722 748 5822 2282
rect 5722 156 5728 748
rect 5816 156 5822 748
rect 5722 0 5822 156
<< via2 >>
rect 971 6539 1089 6657
rect 1247 6539 1365 6657
rect 1523 6539 1641 6657
rect 1799 6539 1917 6657
rect 2075 6539 2193 6657
rect 2351 6539 2469 6657
rect 2627 6539 2745 6657
rect 2903 6539 3021 6657
rect 3179 6539 3297 6657
rect 3455 6539 3573 6657
rect 3731 6539 3849 6657
rect 4007 6539 4125 6657
rect 4283 6539 4401 6657
rect 4559 6539 4677 6657
rect 4835 6539 4953 6657
rect 5111 6539 5229 6657
rect 893 5917 963 5987
rect 1169 5917 1239 5987
rect 1445 5917 1515 5987
rect 1721 5917 1791 5987
rect 1997 5917 2067 5987
rect 2273 5917 2343 5987
rect 2549 5917 2619 5987
rect 2825 5917 2895 5987
rect 3101 5917 3171 5987
rect 3377 5917 3447 5987
rect 3653 5917 3723 5987
rect 3929 5917 3999 5987
rect 4205 5917 4275 5987
rect 4481 5917 4551 5987
rect 4757 5917 4827 5987
rect 5033 5917 5103 5987
rect 4458 5088 4518 5148
rect 4624 5088 4684 5148
rect 4790 5088 4850 5148
rect 4956 5088 5016 5148
rect 5122 5088 5182 5148
rect 5288 5088 5348 5148
rect 4292 5007 4352 5067
rect 4126 4877 4186 4937
rect 3960 4747 4020 4807
rect 155 3317 215 3377
rect 3794 4617 3854 4677
rect 3628 4487 3688 4547
rect 3462 4357 3522 4417
rect 3296 4227 3356 4287
rect 3130 4097 3190 4157
rect 2964 3967 3024 4027
rect 2959 3447 3029 3517
rect 2881 3317 2941 3377
rect 2798 3187 2858 3247
rect 2632 3057 2692 3117
rect 2466 2927 2526 2987
rect 2300 2797 2360 2857
rect 2134 2667 2194 2727
rect 1968 2537 2028 2597
rect 5454 2502 5514 2562
rect 1802 2407 1862 2467
rect 1636 2277 1696 2337
rect 1470 2147 1530 2207
rect 308 2066 368 2126
rect 474 2066 534 2126
rect 640 2066 700 2126
rect 806 2066 866 2126
rect 972 2066 1032 2126
rect 1138 2066 1198 2126
rect 1304 2066 1364 2126
rect 719 1227 789 1297
rect 995 1227 1065 1297
rect 1271 1227 1341 1297
rect 1547 1227 1617 1297
rect 1823 1227 1893 1297
rect 2099 1227 2169 1297
rect 2375 1227 2445 1297
rect 2651 1227 2721 1297
rect 2927 1227 2997 1297
rect 3203 1227 3273 1297
rect 3479 1227 3549 1297
rect 3755 1227 3825 1297
rect 4031 1227 4101 1297
rect 4307 1227 4377 1297
rect 4583 1227 4653 1297
rect 4859 1227 4929 1297
rect 5135 1227 5205 1297
rect 593 557 711 675
rect 869 557 987 675
rect 1145 557 1263 675
rect 1421 557 1539 675
rect 1697 557 1815 675
rect 1973 557 2091 675
rect 2249 557 2367 675
rect 2525 557 2643 675
rect 2801 557 2919 675
rect 3077 557 3195 675
rect 3353 557 3471 675
rect 3629 557 3747 675
rect 3905 557 4023 675
rect 4181 557 4299 675
rect 4457 557 4575 675
rect 4733 557 4851 675
rect 5009 557 5127 675
<< metal3 >>
rect 961 6657 5239 6667
rect 961 6539 971 6657
rect 1089 6539 1247 6657
rect 1365 6539 1523 6657
rect 1641 6539 1799 6657
rect 1917 6539 2075 6657
rect 2193 6539 2351 6657
rect 2469 6539 2627 6657
rect 2745 6539 2903 6657
rect 3021 6539 3179 6657
rect 3297 6539 3455 6657
rect 3573 6539 3731 6657
rect 3849 6539 4007 6657
rect 4125 6539 4283 6657
rect 4401 6539 4559 6657
rect 4677 6539 4835 6657
rect 4953 6539 5111 6657
rect 5229 6539 5239 6657
rect 961 6529 5239 6539
rect 888 5987 968 5992
rect 888 5917 893 5987
rect 963 5917 968 5987
rect 888 5912 968 5917
rect 1164 5987 1244 5992
rect 1164 5917 1169 5987
rect 1239 5917 1244 5987
rect 1164 5912 1244 5917
rect 1440 5987 1520 5992
rect 1440 5917 1445 5987
rect 1515 5917 1520 5987
rect 1440 5912 1520 5917
rect 1716 5987 1796 5992
rect 1716 5917 1721 5987
rect 1791 5917 1796 5987
rect 1716 5912 1796 5917
rect 1992 5987 2072 5992
rect 1992 5917 1997 5987
rect 2067 5917 2072 5987
rect 1992 5912 2072 5917
rect 2268 5987 2348 5992
rect 2268 5917 2273 5987
rect 2343 5917 2348 5987
rect 2268 5912 2348 5917
rect 2544 5987 2624 5992
rect 2544 5917 2549 5987
rect 2619 5917 2624 5987
rect 2544 5912 2624 5917
rect 2820 5987 2900 5992
rect 2820 5917 2825 5987
rect 2895 5917 2900 5987
rect 2820 5912 2900 5917
rect 3096 5987 3176 5992
rect 3096 5917 3101 5987
rect 3171 5917 3176 5987
rect 3096 5912 3176 5917
rect 3372 5987 3452 5992
rect 3372 5917 3377 5987
rect 3447 5917 3452 5987
rect 3372 5912 3452 5917
rect 3648 5987 3728 5992
rect 3648 5917 3653 5987
rect 3723 5917 3728 5987
rect 3648 5912 3728 5917
rect 3924 5987 4004 5992
rect 3924 5917 3929 5987
rect 3999 5917 4004 5987
rect 3924 5912 4004 5917
rect 4200 5987 4280 5992
rect 4200 5917 4205 5987
rect 4275 5917 4280 5987
rect 4200 5912 4280 5917
rect 4476 5987 4556 5992
rect 4476 5917 4481 5987
rect 4551 5917 4556 5987
rect 4476 5912 4556 5917
rect 4752 5987 4832 5992
rect 4752 5917 4757 5987
rect 4827 5917 4832 5987
rect 4752 5912 4832 5917
rect 5028 5987 5108 5992
rect 5028 5917 5033 5987
rect 5103 5917 5519 5987
rect 5028 5912 5108 5917
rect 893 4032 963 5912
rect 1169 4162 1239 5912
rect 1445 4292 1515 5912
rect 1721 4422 1791 5912
rect 1997 4552 2067 5912
rect 2273 4682 2343 5912
rect 2549 4812 2619 5912
rect 2825 4942 2895 5912
rect 3101 5072 3171 5912
rect 3377 5202 3447 5912
rect 3653 5332 3723 5912
rect 3929 5462 3999 5912
rect 4205 5592 4275 5912
rect 4481 5722 4551 5912
rect 4757 5852 4827 5912
rect 4757 5782 5353 5852
rect 4481 5652 5187 5722
rect 4205 5522 5021 5592
rect 3929 5392 4855 5462
rect 3653 5262 4689 5332
rect 3377 5148 4523 5202
rect 3377 5132 4458 5148
rect 4453 5088 4458 5132
rect 4518 5088 4523 5148
rect 4453 5083 4523 5088
rect 4619 5148 4689 5262
rect 4619 5088 4624 5148
rect 4684 5088 4689 5148
rect 4619 5083 4689 5088
rect 4785 5148 4855 5392
rect 4785 5088 4790 5148
rect 4850 5088 4855 5148
rect 4785 5083 4855 5088
rect 4951 5148 5021 5522
rect 4951 5088 4956 5148
rect 5016 5088 5021 5148
rect 4951 5083 5021 5088
rect 5117 5148 5187 5652
rect 5117 5088 5122 5148
rect 5182 5088 5187 5148
rect 5117 5083 5187 5088
rect 5283 5148 5353 5782
rect 5283 5088 5288 5148
rect 5348 5088 5353 5148
rect 5283 5083 5353 5088
rect 3101 5067 4357 5072
rect 3101 5007 4292 5067
rect 4352 5007 4357 5067
rect 3101 5002 4357 5007
rect 2825 4937 4191 4942
rect 2825 4877 4126 4937
rect 4186 4877 4191 4937
rect 2825 4872 4191 4877
rect 2549 4807 4025 4812
rect 2549 4747 3960 4807
rect 4020 4747 4025 4807
rect 2549 4742 4025 4747
rect 2273 4677 3859 4682
rect 2273 4617 3794 4677
rect 3854 4617 3859 4677
rect 2273 4612 3859 4617
rect 1997 4547 3693 4552
rect 1997 4487 3628 4547
rect 3688 4487 3693 4547
rect 1997 4482 3693 4487
rect 1721 4417 3527 4422
rect 1721 4357 3462 4417
rect 3522 4357 3527 4417
rect 1721 4352 3527 4357
rect 1445 4287 3361 4292
rect 1445 4227 3296 4287
rect 3356 4227 3361 4287
rect 1445 4222 3361 4227
rect 1169 4157 3195 4162
rect 1169 4097 3130 4157
rect 3190 4097 3195 4157
rect 1169 4092 3195 4097
rect 893 4027 3029 4032
rect 893 3967 2964 4027
rect 3024 3967 3029 4027
rect 893 3962 3029 3967
rect 2954 3517 3034 3522
rect 2954 3447 2959 3517
rect 3029 3447 5340 3517
rect 2954 3442 3034 3447
rect 150 3377 5205 3382
rect 150 3317 155 3377
rect 215 3317 2881 3377
rect 2941 3317 5205 3377
rect 150 3312 5205 3317
rect 2793 3247 4929 3252
rect 2793 3187 2798 3247
rect 2858 3187 4929 3247
rect 2793 3182 4929 3187
rect 2627 3117 4653 3122
rect 2627 3057 2632 3117
rect 2692 3057 4653 3117
rect 2627 3052 4653 3057
rect 2461 2987 4377 2992
rect 2461 2927 2466 2987
rect 2526 2927 4377 2987
rect 2461 2922 4377 2927
rect 2295 2857 4101 2862
rect 2295 2797 2300 2857
rect 2360 2797 4101 2857
rect 2295 2792 4101 2797
rect 2129 2727 3825 2732
rect 2129 2667 2134 2727
rect 2194 2667 3825 2727
rect 2129 2662 3825 2667
rect 1963 2597 3549 2602
rect 1963 2537 1968 2597
rect 2028 2537 3549 2597
rect 1963 2532 3549 2537
rect 1797 2467 3273 2472
rect 1797 2407 1802 2467
rect 1862 2407 3273 2467
rect 1797 2402 3273 2407
rect 1631 2337 2997 2342
rect 1631 2277 1636 2337
rect 1696 2277 2997 2337
rect 1631 2272 2997 2277
rect 1465 2207 2721 2212
rect 1465 2147 1470 2207
rect 1530 2147 2721 2207
rect 1465 2142 2721 2147
rect 303 2126 373 2131
rect 303 2066 308 2126
rect 368 2066 373 2126
rect 303 1297 373 2066
rect 469 2126 539 2131
rect 469 2066 474 2126
rect 534 2066 539 2126
rect 469 1432 539 2066
rect 635 2126 705 2131
rect 635 2066 640 2126
rect 700 2066 705 2126
rect 635 1562 705 2066
rect 801 2126 871 2131
rect 801 2066 806 2126
rect 866 2066 871 2126
rect 801 1692 871 2066
rect 967 2126 1037 2131
rect 967 2066 972 2126
rect 1032 2066 1037 2126
rect 967 1822 1037 2066
rect 1133 2126 1203 2131
rect 1133 2066 1138 2126
rect 1198 2066 1203 2126
rect 1133 1952 1203 2066
rect 1299 2126 1369 2131
rect 1299 2066 1304 2126
rect 1364 2082 1369 2126
rect 1364 2066 2445 2082
rect 1299 2012 2445 2066
rect 1133 1882 2169 1952
rect 967 1752 1893 1822
rect 801 1622 1617 1692
rect 635 1492 1341 1562
rect 469 1362 1065 1432
rect 995 1302 1065 1362
rect 1271 1302 1341 1492
rect 1547 1302 1617 1622
rect 1823 1302 1893 1752
rect 2099 1302 2169 1882
rect 2375 1302 2445 2012
rect 2651 1302 2721 2142
rect 2927 1302 2997 2272
rect 3203 1302 3273 2402
rect 3479 1302 3549 2532
rect 3755 1302 3825 2662
rect 4031 1302 4101 2792
rect 4307 1302 4377 2922
rect 4583 1302 4653 3052
rect 4859 1302 4929 3182
rect 5135 1302 5205 3312
rect 714 1297 794 1302
rect 303 1227 719 1297
rect 789 1227 794 1297
rect 714 1222 794 1227
rect 990 1297 1070 1302
rect 990 1227 995 1297
rect 1065 1227 1070 1297
rect 990 1222 1070 1227
rect 1266 1297 1346 1302
rect 1266 1227 1271 1297
rect 1341 1227 1346 1297
rect 1266 1222 1346 1227
rect 1542 1297 1622 1302
rect 1542 1227 1547 1297
rect 1617 1227 1622 1297
rect 1542 1222 1622 1227
rect 1818 1297 1898 1302
rect 1818 1227 1823 1297
rect 1893 1227 1898 1297
rect 1818 1222 1898 1227
rect 2094 1297 2174 1302
rect 2094 1227 2099 1297
rect 2169 1227 2174 1297
rect 2094 1222 2174 1227
rect 2370 1297 2450 1302
rect 2370 1227 2375 1297
rect 2445 1227 2450 1297
rect 2370 1222 2450 1227
rect 2646 1297 2726 1302
rect 2646 1227 2651 1297
rect 2721 1227 2726 1297
rect 2646 1222 2726 1227
rect 2922 1297 3002 1302
rect 2922 1227 2927 1297
rect 2997 1227 3002 1297
rect 2922 1222 3002 1227
rect 3198 1297 3278 1302
rect 3198 1227 3203 1297
rect 3273 1227 3278 1297
rect 3198 1222 3278 1227
rect 3474 1297 3554 1302
rect 3474 1227 3479 1297
rect 3549 1227 3554 1297
rect 3474 1222 3554 1227
rect 3750 1297 3830 1302
rect 3750 1227 3755 1297
rect 3825 1227 3830 1297
rect 3750 1222 3830 1227
rect 4026 1297 4106 1302
rect 4026 1227 4031 1297
rect 4101 1227 4106 1297
rect 4026 1222 4106 1227
rect 4302 1297 4382 1302
rect 4302 1227 4307 1297
rect 4377 1227 4382 1297
rect 4302 1222 4382 1227
rect 4578 1297 4658 1302
rect 4578 1227 4583 1297
rect 4653 1227 4658 1297
rect 4578 1222 4658 1227
rect 4854 1297 4934 1302
rect 4854 1227 4859 1297
rect 4929 1227 4934 1297
rect 4854 1222 4934 1227
rect 5130 1297 5210 1302
rect 5130 1227 5135 1297
rect 5205 1227 5210 1297
rect 5130 1222 5210 1227
rect 5270 815 5340 3447
rect 5449 2572 5519 5917
rect 5444 2562 5524 2572
rect 5444 2502 5454 2562
rect 5514 2502 5524 2562
rect 5444 2492 5524 2502
rect 893 745 5340 815
rect 893 685 963 745
rect 1445 685 1515 745
rect 1997 685 2067 745
rect 2549 685 2619 745
rect 3101 685 3171 745
rect 3653 685 3723 745
rect 4205 685 4275 745
rect 4757 685 4827 745
rect 583 675 721 685
rect 583 557 593 675
rect 711 557 721 675
rect 583 547 721 557
rect 859 675 997 685
rect 859 557 869 675
rect 987 557 997 675
rect 859 547 997 557
rect 1135 675 1273 685
rect 1135 557 1145 675
rect 1263 557 1273 675
rect 1135 547 1273 557
rect 1411 675 1549 685
rect 1411 557 1421 675
rect 1539 557 1549 675
rect 1411 547 1549 557
rect 1687 675 1825 685
rect 1687 557 1697 675
rect 1815 557 1825 675
rect 1687 547 1825 557
rect 1963 675 2101 685
rect 1963 557 1973 675
rect 2091 557 2101 675
rect 1963 547 2101 557
rect 2239 675 2377 685
rect 2239 557 2249 675
rect 2367 557 2377 675
rect 2239 547 2377 557
rect 2515 675 2653 685
rect 2515 557 2525 675
rect 2643 557 2653 675
rect 2515 547 2653 557
rect 2791 675 2929 685
rect 2791 557 2801 675
rect 2919 557 2929 675
rect 2791 547 2929 557
rect 3067 675 3205 685
rect 3067 557 3077 675
rect 3195 557 3205 675
rect 3067 547 3205 557
rect 3343 675 3481 685
rect 3343 557 3353 675
rect 3471 557 3481 675
rect 3343 547 3481 557
rect 3619 675 3757 685
rect 3619 557 3629 675
rect 3747 557 3757 675
rect 3619 547 3757 557
rect 3895 675 4033 685
rect 3895 557 3905 675
rect 4023 557 4033 675
rect 3895 547 4033 557
rect 4171 675 4309 685
rect 4171 557 4181 675
rect 4299 557 4309 675
rect 4171 547 4309 557
rect 4447 675 4585 685
rect 4447 557 4457 675
rect 4575 557 4585 675
rect 4447 547 4585 557
rect 4723 675 4861 685
rect 4723 557 4733 675
rect 4851 557 4861 675
rect 4723 547 4861 557
rect 4999 675 5137 685
rect 4999 557 5009 675
rect 5127 557 5137 675
rect 4999 547 5137 557
rect 617 487 687 547
rect 1169 487 1239 547
rect 1721 487 1791 547
rect 2273 487 2343 547
rect 2825 487 2895 547
rect 3377 487 3447 547
rect 3929 487 3999 547
rect 4481 487 4551 547
rect 5033 487 5103 547
rect 5449 487 5519 2492
rect 617 417 5519 487
use passgates  passgates_0
timestamp 1740604869
transform -1 0 5681 0 -1 7214
box 0 0 5540 2076
use passgates  passgates_2
timestamp 1740604869
transform 1 0 141 0 1 0
box 0 0 5540 2076
use sky130_fd_pr__res_xhigh_po_0p35_7C4M5Y  sky130_fd_pr__res_xhigh_po_0p35_7C4M5Y_0
timestamp 1740618740
transform 1 0 2911 0 1 3607
box -2911 -1511 2911 1511
<< labels >>
flabel metal2 0 0 100 7214 1 FreeSans 400 0 0 0 VSS
port 1 n ground bidirectional
flabel metal2 150 0 250 7214 1 FreeSans 400 0 0 0 VDD
port 2 n power bidirectional
flabel metal3 961 6529 5239 6667 1 FreeSans 400 0 0 0 VOUT
port 3 n signal default
flabel metal3 617 417 5519 487 1 FreeSans 400 0 0 0 A
flabel metal3 893 745 5340 815 1 FreeSans 400 0 0 0 B
flabel metal2 5101 6701 5239 6839 1 FreeSans 400 0 0 0 D[0]
port 4 n signal default
flabel metal2 4825 6701 4963 6839 1 FreeSans 400 0 0 0 D[1]
port 5 n signal default
flabel metal2 4549 6701 4687 6839 1 FreeSans 400 0 0 0 D[2]
port 6 n signal default
flabel metal2 4273 6701 4411 6839 1 FreeSans 400 0 0 0 D[3]
port 7 n signal default
flabel metal2 3997 6701 4135 6839 1 FreeSans 400 0 0 0 D[4]
port 8 n signal default
flabel metal2 3721 6701 3859 6839 1 FreeSans 400 0 0 0 D[5]
port 9 n signal default
flabel metal2 3445 6701 3583 6839 1 FreeSans 400 0 0 0 D[6]
port 10 n signal default
flabel metal2 3169 6701 3307 6839 1 FreeSans 400 0 0 0 D[7]
port 11 n signal default
flabel metal2 2893 6701 3031 6839 1 FreeSans 400 0 0 0 D[8]
port 12 n signal default
flabel metal2 2617 6701 2755 6839 1 FreeSans 400 0 0 0 D[9]
port 13 n signal default
flabel metal2 2341 6701 2479 6839 1 FreeSans 400 0 0 0 D[10]
port 14 n signal default
flabel metal2 2065 6701 2203 6839 1 FreeSans 400 0 0 0 D[11]
port 15 n signal default
flabel metal2 1789 6701 1927 6839 1 FreeSans 400 0 0 0 D[12]
port 16 n signal default
flabel metal2 1513 6701 1651 6839 1 FreeSans 400 0 0 0 D[13]
port 17 n signal default
flabel metal2 1237 6701 1375 6839 1 FreeSans 400 0 0 0 D[14]
port 18 n signal default
flabel metal2 961 6701 1099 6839 1 FreeSans 400 0 0 0 D[15]
port 19 n signal default
flabel metal2 583 375 721 513 1 FreeSans 400 0 0 0 C[0]
port 20 n signal default
flabel metal2 859 375 997 513 1 FreeSans 400 0 0 0 C[1]
port 21 n signal default
flabel metal2 1135 375 1273 513 1 FreeSans 400 0 0 0 C[2]
port 22 n signal default
flabel metal2 1411 375 1549 513 1 FreeSans 400 0 0 0 C[3]
port 23 n signal default
flabel metal2 1687 375 1825 513 1 FreeSans 400 0 0 0 C[4]
port 24 n signal default
flabel metal2 1963 375 2101 513 1 FreeSans 400 0 0 0 C[5]
port 25 n signal default
flabel metal2 2239 375 2377 513 1 FreeSans 400 0 0 0 C[6]
port 26 n signal default
flabel metal2 2515 375 2653 513 1 FreeSans 400 0 0 0 C[7]
port 27 n signal default
flabel metal2 2791 375 2929 513 1 FreeSans 400 0 0 0 C[8]
port 28 n signal default
flabel metal2 3067 375 3205 513 1 FreeSans 400 0 0 0 C[9]
port 29 n signal default
flabel metal2 3343 375 3481 513 1 FreeSans 400 0 0 0 C[10]
port 30 n signal default
flabel metal2 3619 375 3757 513 1 FreeSans 400 0 0 0 C[11]
port 31 n signal default
flabel metal2 3895 375 4033 513 1 FreeSans 400 0 0 0 C[12]
port 32 n signal default
flabel metal2 4171 375 4309 513 1 FreeSans 400 0 0 0 C[13]
port 33 n signal default
flabel metal2 4447 375 4585 513 1 FreeSans 400 0 0 0 C[14]
port 34 n signal default
flabel metal2 4723 375 4861 513 1 FreeSans 400 0 0 0 C[15]
port 35 n signal default
flabel metal2 4999 375 5137 513 1 FreeSans 400 0 0 0 C[16]
port 36 n signal default
<< end >>
