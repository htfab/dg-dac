magic
tech sky130A
magscale 1 2
timestamp 1748333863
<< metal1 >>
rect 4807 20376 4813 20428
rect 4865 20376 4871 20428
rect 7503 20376 7509 20428
rect 7561 20376 7567 20428
rect 10199 20376 10205 20428
rect 10257 20376 10263 20428
rect 12595 20382 12601 20434
rect 12653 20382 12659 20434
rect 12895 20376 12901 20428
rect 12953 20376 12959 20428
rect 5899 15860 5951 15866
rect 13776 15860 13828 15866
rect 5951 15817 13776 15851
rect 5899 15802 5951 15808
rect 13776 15802 13828 15808
rect 6175 15783 6227 15789
rect 14473 15783 14525 15789
rect 6227 15740 14473 15774
rect 6175 15725 6227 15731
rect 14473 15725 14525 15731
rect 6451 15706 6503 15712
rect 12434 15706 12486 15712
rect 6503 15663 12434 15697
rect 6451 15648 6503 15654
rect 12434 15648 12486 15654
rect 6727 15629 6779 15635
rect 13131 15629 13183 15635
rect 6779 15586 13131 15620
rect 6727 15571 6779 15577
rect 13131 15571 13183 15577
rect 7003 15552 7055 15558
rect 11092 15552 11144 15558
rect 7055 15509 11092 15543
rect 7003 15494 7055 15500
rect 11092 15494 11144 15500
rect 7279 15475 7331 15481
rect 11789 15475 11841 15481
rect 7331 15432 11789 15466
rect 7279 15417 7331 15423
rect 11789 15417 11841 15423
rect 7555 15398 7607 15404
rect 9750 15398 9802 15404
rect 7607 15355 9750 15389
rect 7555 15340 7607 15346
rect 9750 15340 9802 15346
rect 7831 15321 7883 15327
rect 10447 15321 10499 15327
rect 7883 15278 10447 15312
rect 7831 15263 7883 15269
rect 10447 15263 10499 15269
rect 8107 15244 8159 15250
rect 8482 15244 8534 15250
rect 8159 15201 8482 15235
rect 8107 15186 8159 15192
rect 8482 15186 8534 15192
rect 8383 15167 8435 15173
rect 9105 15167 9157 15173
rect 8435 15124 9105 15158
rect 8383 15109 8435 15115
rect 9105 15109 9157 15115
rect 7140 15090 7192 15096
rect 8659 15090 8711 15096
rect 7192 15047 8659 15081
rect 7140 15032 7192 15038
rect 8659 15032 8711 15038
rect 7689 15013 7741 15019
rect 8935 15013 8987 15019
rect 7741 14970 8935 15004
rect 7689 14955 7741 14961
rect 8935 14955 8987 14961
rect 4382 14936 4434 14942
rect 5724 14936 5776 14942
rect 4434 14893 5510 14927
rect 4382 14878 4434 14884
rect 5079 14859 5131 14865
rect 5131 14816 5433 14850
rect 5079 14801 5131 14807
rect 5399 14696 5433 14816
rect 5476 14773 5510 14893
rect 9211 14936 9263 14942
rect 5776 14893 9211 14927
rect 5724 14878 5776 14884
rect 9211 14878 9263 14884
rect 6347 14859 6399 14865
rect 9487 14859 9539 14865
rect 6399 14816 9487 14850
rect 6347 14801 6399 14807
rect 9487 14801 9539 14807
rect 9763 14782 9815 14788
rect 5476 14739 9763 14773
rect 9763 14724 9815 14730
rect 10039 14705 10091 14711
rect 5399 14662 10039 14696
rect 10039 14647 10091 14653
rect 7729 6940 7781 6946
rect 8163 6940 8215 6946
rect 7781 6897 8163 6931
rect 7729 6882 7781 6888
rect 8163 6882 8215 6888
rect 963 6863 1015 6869
rect 5521 6863 5573 6869
rect 1015 6820 5521 6854
rect 963 6805 1015 6811
rect 5521 6805 5573 6811
rect 8005 6863 8057 6869
rect 8986 6863 9038 6869
rect 8057 6820 8986 6854
rect 8005 6805 8057 6811
rect 8986 6805 9038 6811
rect 1863 6786 1915 6792
rect 5797 6786 5849 6792
rect 1915 6743 5797 6777
rect 1863 6728 1915 6734
rect 5797 6728 5849 6734
rect 8281 6786 8333 6792
rect 10040 6786 10092 6792
rect 8333 6743 10040 6777
rect 8281 6728 8333 6734
rect 10040 6728 10092 6734
rect 2763 6709 2815 6715
rect 6073 6709 6125 6715
rect 2815 6666 6073 6700
rect 2763 6651 2815 6657
rect 6073 6651 6125 6657
rect 8557 6709 8609 6715
rect 10863 6709 10915 6715
rect 8609 6666 10863 6700
rect 8557 6651 8609 6657
rect 10863 6651 10915 6657
rect 3663 6632 3715 6638
rect 6349 6632 6401 6638
rect 3715 6589 6349 6623
rect 3663 6574 3715 6580
rect 6349 6574 6401 6580
rect 8833 6632 8885 6638
rect 11763 6632 11815 6638
rect 8885 6589 11763 6623
rect 8833 6574 8885 6580
rect 11763 6574 11815 6580
rect 4563 6555 4615 6561
rect 6625 6555 6677 6561
rect 4615 6512 6625 6546
rect 4563 6497 4615 6503
rect 6625 6497 6677 6503
rect 9109 6555 9161 6561
rect 12663 6555 12715 6561
rect 9161 6512 12663 6546
rect 9109 6497 9161 6503
rect 12663 6497 12715 6503
rect 5463 6478 5515 6484
rect 6901 6478 6953 6484
rect 5515 6435 6901 6469
rect 5463 6420 5515 6426
rect 6901 6420 6953 6426
rect 9385 6478 9437 6484
rect 13563 6478 13615 6484
rect 9437 6435 13563 6469
rect 9385 6420 9437 6426
rect 13563 6420 13615 6426
rect 6363 6401 6415 6407
rect 7177 6401 7229 6407
rect 6415 6358 7177 6392
rect 6363 6343 6415 6349
rect 7177 6343 7229 6349
rect 9661 6401 9713 6407
rect 14463 6401 14515 6407
rect 9713 6358 14463 6392
rect 9661 6343 9713 6349
rect 14463 6343 14515 6349
rect 7263 6324 7315 6330
rect 7453 6324 7505 6330
rect 7315 6281 7453 6315
rect 7263 6266 7315 6272
rect 7453 6266 7505 6272
rect 9937 6324 9989 6330
rect 15363 6324 15415 6330
rect 9989 6281 15363 6315
rect 9937 6266 9989 6272
rect 15363 6266 15415 6272
rect 963 6038 1015 6044
rect 963 5980 1015 5986
rect 1863 6038 1915 6044
rect 1863 5980 1915 5986
rect 2763 6038 2815 6044
rect 2763 5980 2815 5986
rect 3663 6038 3715 6044
rect 3663 5980 3715 5986
rect 4563 6038 4615 6044
rect 4563 5980 4615 5986
rect 5463 6038 5515 6044
rect 5463 5980 5515 5986
rect 6363 6038 6415 6044
rect 6363 5980 6415 5986
rect 7263 6038 7315 6044
rect 7263 5980 7315 5986
rect 8163 6038 8215 6044
rect 8163 5980 8215 5986
rect 9063 6038 9115 6044
rect 9063 5980 9115 5986
rect 9963 6038 10015 6044
rect 9963 5980 10015 5986
rect 10863 6038 10915 6044
rect 10863 5980 10915 5986
rect 11763 6038 11815 6044
rect 11763 5980 11815 5986
rect 12663 6038 12715 6044
rect 12663 5980 12715 5986
rect 13563 6038 13615 6044
rect 13563 5980 13615 5986
rect 14463 6038 14515 6044
rect 14463 5980 14515 5986
rect 15363 6038 15415 6044
rect 15363 5980 15415 5986
<< via1 >>
rect 4813 20376 4865 20428
rect 7509 20376 7561 20428
rect 10205 20376 10257 20428
rect 12601 20382 12653 20434
rect 12901 20376 12953 20428
rect 5899 15808 5951 15860
rect 13776 15808 13828 15860
rect 6175 15731 6227 15783
rect 14473 15731 14525 15783
rect 6451 15654 6503 15706
rect 12434 15654 12486 15706
rect 6727 15577 6779 15629
rect 13131 15577 13183 15629
rect 7003 15500 7055 15552
rect 11092 15500 11144 15552
rect 7279 15423 7331 15475
rect 11789 15423 11841 15475
rect 7555 15346 7607 15398
rect 9750 15346 9802 15398
rect 7831 15269 7883 15321
rect 10447 15269 10499 15321
rect 8107 15192 8159 15244
rect 8482 15192 8534 15244
rect 8383 15115 8435 15167
rect 9105 15115 9157 15167
rect 7140 15038 7192 15090
rect 8659 15038 8711 15090
rect 7689 14961 7741 15013
rect 8935 14961 8987 15013
rect 4382 14884 4434 14936
rect 5079 14807 5131 14859
rect 5724 14884 5776 14936
rect 9211 14884 9263 14936
rect 6347 14807 6399 14859
rect 9487 14807 9539 14859
rect 9763 14730 9815 14782
rect 10039 14653 10091 14705
rect 7729 6888 7781 6940
rect 8163 6888 8215 6940
rect 963 6811 1015 6863
rect 5521 6811 5573 6863
rect 8005 6811 8057 6863
rect 8986 6811 9038 6863
rect 1863 6734 1915 6786
rect 5797 6734 5849 6786
rect 8281 6734 8333 6786
rect 10040 6734 10092 6786
rect 2763 6657 2815 6709
rect 6073 6657 6125 6709
rect 8557 6657 8609 6709
rect 10863 6657 10915 6709
rect 3663 6580 3715 6632
rect 6349 6580 6401 6632
rect 8833 6580 8885 6632
rect 11763 6580 11815 6632
rect 4563 6503 4615 6555
rect 6625 6503 6677 6555
rect 9109 6503 9161 6555
rect 12663 6503 12715 6555
rect 5463 6426 5515 6478
rect 6901 6426 6953 6478
rect 9385 6426 9437 6478
rect 13563 6426 13615 6478
rect 6363 6349 6415 6401
rect 7177 6349 7229 6401
rect 9661 6349 9713 6401
rect 14463 6349 14515 6401
rect 7263 6272 7315 6324
rect 7453 6272 7505 6324
rect 9937 6272 9989 6324
rect 15363 6272 15415 6324
rect 963 5986 1015 6038
rect 1863 5986 1915 6038
rect 2763 5986 2815 6038
rect 3663 5986 3715 6038
rect 4563 5986 4615 6038
rect 5463 5986 5515 6038
rect 6363 5986 6415 6038
rect 7263 5986 7315 6038
rect 8163 5986 8215 6038
rect 9063 5986 9115 6038
rect 9963 5986 10015 6038
rect 10863 5986 10915 6038
rect 11763 5986 11815 6038
rect 12663 5986 12715 6038
rect 13563 5986 13615 6038
rect 14463 5986 14515 6038
rect 15363 5986 15415 6038
<< metal2 >>
rect 16632 21033 16688 21042
rect 4822 20988 16632 21022
rect 490 19785 499 19975
rect 689 19785 698 19975
rect 564 18653 624 19785
rect 864 19575 924 20465
rect 4822 20434 4856 20988
rect 16632 20968 16688 20977
rect 16506 20951 16562 20960
rect 7518 20906 16506 20940
rect 7518 20434 7552 20906
rect 16506 20886 16562 20895
rect 16884 20869 16940 20878
rect 10214 20824 16884 20858
rect 10214 20434 10248 20824
rect 16884 20804 16940 20813
rect 16380 20787 16436 20796
rect 12610 20742 16380 20776
rect 12610 20440 12644 20742
rect 16380 20722 16436 20731
rect 16758 20705 16814 20714
rect 12910 20660 16758 20694
rect 12601 20434 12653 20440
rect 12910 20434 12944 20660
rect 16758 20640 16814 20649
rect 4813 20428 4865 20434
rect 4813 20370 4865 20376
rect 7509 20428 7561 20434
rect 7509 20370 7561 20376
rect 10205 20428 10257 20434
rect 12601 20376 12653 20382
rect 12901 20428 12953 20434
rect 10205 20370 10257 20376
rect 12901 20370 12953 20376
rect 14672 19575 14732 20465
rect 14898 19785 14907 19975
rect 15097 19785 15106 19975
rect 790 19385 799 19575
rect 989 19385 998 19575
rect 14599 19385 14608 19575
rect 14798 19385 14807 19575
rect 864 18353 924 19385
rect 14672 18353 14732 19385
rect 14972 18653 15032 19785
rect 564 15575 624 16797
rect 488 15385 497 15575
rect 687 15385 696 15575
rect 864 15175 924 17097
rect 790 14985 799 15175
rect 989 14985 998 15175
rect 4391 14936 4425 15980
rect 4769 14985 4778 15175
rect 4968 14985 4977 15175
rect 4376 14884 4382 14936
rect 4434 14884 4440 14936
rect 4823 14684 4923 14985
rect 5088 14859 5122 15980
rect 5273 15385 5282 15575
rect 5472 15385 5481 15575
rect 5073 14807 5079 14859
rect 5131 14807 5137 14859
rect 5327 14684 5427 15385
rect 5733 14936 5767 15980
rect 5893 15808 5899 15860
rect 5951 15808 5957 15860
rect 5718 14884 5724 14936
rect 5776 14884 5782 14936
rect 4823 14584 4995 14684
rect 4895 14382 4995 14584
rect 5045 14584 5427 14684
rect 5045 14382 5145 14584
rect 5908 14570 5942 15808
rect 6169 15731 6175 15783
rect 6227 15731 6233 15783
rect 6430 15774 6464 15980
rect 6356 15740 6464 15774
rect 6184 14570 6218 15731
rect 6356 14859 6390 15740
rect 6445 15654 6451 15706
rect 6503 15654 6509 15706
rect 6341 14807 6347 14859
rect 6399 14807 6405 14859
rect 6460 14570 6494 15654
rect 6721 15577 6727 15629
rect 6779 15577 6785 15629
rect 7075 15620 7109 15980
rect 7075 15586 7183 15620
rect 6736 14570 6770 15577
rect 6997 15500 7003 15552
rect 7055 15500 7061 15552
rect 7012 14570 7046 15500
rect 7149 15090 7183 15586
rect 7273 15423 7279 15475
rect 7331 15423 7337 15475
rect 7134 15038 7140 15090
rect 7192 15038 7198 15090
rect 7288 14570 7322 15423
rect 7549 15346 7555 15398
rect 7607 15346 7613 15398
rect 7772 15389 7806 15980
rect 7698 15355 7806 15389
rect 7564 14570 7598 15346
rect 7698 15013 7732 15355
rect 7825 15269 7831 15321
rect 7883 15269 7889 15321
rect 8417 15312 8451 15980
rect 8417 15278 8525 15312
rect 7683 14961 7689 15013
rect 7741 14961 7747 15013
rect 7840 14570 7874 15269
rect 8491 15244 8525 15278
rect 8101 15192 8107 15244
rect 8159 15192 8165 15244
rect 8476 15192 8482 15244
rect 8534 15192 8540 15244
rect 8116 14570 8150 15192
rect 9114 15167 9148 15980
rect 9759 15398 9793 15980
rect 9744 15346 9750 15398
rect 9802 15346 9808 15398
rect 10164 15385 10173 15575
rect 10363 15385 10372 15575
rect 8377 15115 8383 15167
rect 8435 15115 8441 15167
rect 9099 15115 9105 15167
rect 9157 15115 9163 15167
rect 8392 14570 8426 15115
rect 8653 15038 8659 15090
rect 8711 15038 8717 15090
rect 8668 14570 8702 15038
rect 8929 14961 8935 15013
rect 8987 14961 8993 15013
rect 8944 14570 8978 14961
rect 9205 14884 9211 14936
rect 9263 14884 9269 14936
rect 10218 14884 10318 15385
rect 10456 15321 10490 15980
rect 11101 15552 11135 15980
rect 11086 15500 11092 15552
rect 11144 15500 11150 15552
rect 11798 15475 11832 15980
rect 12443 15706 12477 15980
rect 12428 15654 12434 15706
rect 12486 15654 12492 15706
rect 13140 15629 13174 15980
rect 13785 15860 13819 15980
rect 13770 15808 13776 15860
rect 13828 15808 13834 15860
rect 14482 15783 14516 15980
rect 14467 15731 14473 15783
rect 14525 15731 14531 15783
rect 13125 15577 13131 15629
rect 13183 15577 13189 15629
rect 11783 15423 11789 15475
rect 11841 15423 11847 15475
rect 10441 15269 10447 15321
rect 10499 15269 10505 15321
rect 14672 15175 14732 17097
rect 14972 15575 15032 16797
rect 14897 15385 14906 15575
rect 15096 15385 15105 15575
rect 10565 14985 10574 15175
rect 10764 14985 10773 15175
rect 14599 14985 14608 15175
rect 14798 14985 14807 15175
rect 9220 14570 9254 14884
rect 9481 14807 9487 14859
rect 9539 14807 9545 14859
rect 9496 14570 9530 14807
rect 10218 14784 10567 14884
rect 9757 14730 9763 14782
rect 9815 14730 9821 14782
rect 9772 14570 9806 14730
rect 10033 14653 10039 14705
rect 10091 14653 10097 14705
rect 10048 14570 10082 14653
rect 5888 14514 5897 14570
rect 5953 14514 5962 14570
rect 6164 14514 6173 14570
rect 6229 14514 6238 14570
rect 6440 14514 6449 14570
rect 6505 14514 6514 14570
rect 6716 14514 6725 14570
rect 6781 14514 6790 14570
rect 6992 14514 7001 14570
rect 7057 14514 7066 14570
rect 7268 14514 7277 14570
rect 7333 14514 7342 14570
rect 7544 14514 7553 14570
rect 7609 14514 7618 14570
rect 7820 14514 7829 14570
rect 7885 14514 7894 14570
rect 8096 14514 8105 14570
rect 8161 14514 8170 14570
rect 8372 14514 8381 14570
rect 8437 14514 8446 14570
rect 8648 14514 8657 14570
rect 8713 14514 8722 14570
rect 8924 14514 8933 14570
rect 8989 14514 8998 14570
rect 9200 14514 9209 14570
rect 9265 14514 9274 14570
rect 9476 14514 9485 14570
rect 9541 14514 9550 14570
rect 9752 14514 9761 14570
rect 9817 14514 9826 14570
rect 10028 14514 10037 14570
rect 10093 14514 10102 14570
rect 10467 14382 10567 14784
rect 10617 14382 10717 14985
rect 5895 14235 5955 14244
rect 5895 14008 5955 14179
rect 6171 14235 6231 14244
rect 6171 14008 6231 14179
rect 6447 14235 6507 14244
rect 6447 14008 6507 14179
rect 6723 14235 6783 14244
rect 6723 14008 6783 14179
rect 6999 14235 7059 14244
rect 6999 14008 7059 14179
rect 7275 14235 7335 14244
rect 7275 14008 7335 14179
rect 7551 14235 7611 14244
rect 7551 14008 7611 14179
rect 7827 14235 7887 14244
rect 7827 14008 7887 14179
rect 8103 14235 8163 14244
rect 8103 14008 8163 14179
rect 8379 14235 8439 14244
rect 8379 14008 8439 14179
rect 8655 14235 8715 14244
rect 8655 14008 8715 14179
rect 8931 14235 8991 14244
rect 8931 14008 8991 14179
rect 9207 14235 9267 14244
rect 9207 14008 9267 14179
rect 9483 14235 9543 14244
rect 9483 14008 9543 14179
rect 9759 14235 9819 14244
rect 9759 14008 9819 14179
rect 10035 14235 10095 14244
rect 10035 14008 10095 14179
rect 5517 7393 5577 7562
rect 5517 7328 5577 7337
rect 5793 7393 5853 7562
rect 5793 7328 5853 7337
rect 6069 7393 6129 7562
rect 6069 7328 6129 7337
rect 6345 7393 6405 7562
rect 6345 7328 6405 7337
rect 6621 7393 6681 7562
rect 6621 7328 6681 7337
rect 6897 7393 6957 7562
rect 6897 7328 6957 7337
rect 7173 7393 7233 7562
rect 7173 7328 7233 7337
rect 7449 7393 7509 7562
rect 7449 7328 7509 7337
rect 7725 7393 7785 7562
rect 7725 7328 7785 7337
rect 8001 7393 8061 7562
rect 8001 7328 8061 7337
rect 8277 7393 8337 7562
rect 8277 7328 8337 7337
rect 8553 7393 8613 7562
rect 8553 7328 8613 7337
rect 8829 7393 8889 7562
rect 8829 7328 8889 7337
rect 9105 7393 9165 7562
rect 9105 7328 9165 7337
rect 9381 7393 9441 7562
rect 9381 7328 9441 7337
rect 9657 7393 9717 7562
rect 9657 7328 9717 7337
rect 9933 7393 9993 7562
rect 9933 7328 9993 7337
rect 4840 7088 4995 7188
rect 957 6811 963 6863
rect 1015 6811 1021 6863
rect -4 6405 5 6595
rect 195 6405 204 6595
rect 65 4432 125 6405
rect 972 6038 1006 6811
rect 1857 6734 1863 6786
rect 1915 6734 1921 6786
rect 957 5986 963 6038
rect 1015 5986 1021 6038
rect 1204 6005 1213 6195
rect 1403 6005 1412 6195
rect 1872 6038 1906 6734
rect 2757 6657 2763 6709
rect 2815 6657 2821 6709
rect 2772 6038 2806 6657
rect 3657 6580 3663 6632
rect 3715 6580 3721 6632
rect 3672 6038 3706 6580
rect 4557 6503 4563 6555
rect 4615 6503 4621 6555
rect 4572 6038 4606 6503
rect 4840 6195 4940 7088
rect 5045 6595 5145 7188
rect 5510 7004 5519 7060
rect 5575 7004 5584 7060
rect 5786 7004 5795 7060
rect 5851 7004 5860 7060
rect 6062 7004 6071 7060
rect 6127 7004 6136 7060
rect 6338 7004 6347 7060
rect 6403 7004 6412 7060
rect 6614 7004 6623 7060
rect 6679 7004 6688 7060
rect 6890 7004 6899 7060
rect 6955 7004 6964 7060
rect 7166 7004 7175 7060
rect 7231 7004 7240 7060
rect 7442 7004 7451 7060
rect 7507 7004 7516 7060
rect 7718 7004 7727 7060
rect 7783 7004 7792 7060
rect 7994 7004 8003 7060
rect 8059 7004 8068 7060
rect 8270 7004 8279 7060
rect 8335 7004 8344 7060
rect 8546 7004 8555 7060
rect 8611 7004 8620 7060
rect 8822 7004 8831 7060
rect 8887 7004 8896 7060
rect 9098 7004 9107 7060
rect 9163 7004 9172 7060
rect 9374 7004 9383 7060
rect 9439 7004 9448 7060
rect 9650 7004 9659 7060
rect 9715 7004 9724 7060
rect 9926 7004 9935 7060
rect 9991 7004 10000 7060
rect 5530 6863 5564 7004
rect 5515 6811 5521 6863
rect 5573 6811 5579 6863
rect 5806 6786 5840 7004
rect 5791 6734 5797 6786
rect 5849 6734 5855 6786
rect 6082 6709 6116 7004
rect 6067 6657 6073 6709
rect 6125 6657 6131 6709
rect 6358 6632 6392 7004
rect 4989 6405 4998 6595
rect 5188 6405 5197 6595
rect 6343 6580 6349 6632
rect 6401 6580 6407 6632
rect 6634 6555 6668 7004
rect 6619 6503 6625 6555
rect 6677 6503 6683 6555
rect 6910 6478 6944 7004
rect 5457 6426 5463 6478
rect 5515 6426 5521 6478
rect 6895 6426 6901 6478
rect 6953 6426 6959 6478
rect 1278 5815 1338 6005
rect 1857 5986 1863 6038
rect 1915 5986 1921 6038
rect 2757 5986 2763 6038
rect 2815 5986 2821 6038
rect 3657 5986 3663 6038
rect 3715 5986 3721 6038
rect 4557 5986 4563 6038
rect 4615 5986 4621 6038
rect 4786 6005 4795 6195
rect 4985 6005 4994 6195
rect 5472 6038 5506 6426
rect 7186 6401 7220 7004
rect 6357 6349 6363 6401
rect 6415 6349 6421 6401
rect 7171 6349 7177 6401
rect 7229 6349 7235 6401
rect 6372 6038 6406 6349
rect 7462 6324 7496 7004
rect 7738 6940 7772 7004
rect 7723 6888 7729 6940
rect 7781 6888 7787 6940
rect 8014 6863 8048 7004
rect 8157 6888 8163 6940
rect 8215 6888 8221 6940
rect 7999 6811 8005 6863
rect 8057 6811 8063 6863
rect 7257 6272 7263 6324
rect 7315 6272 7321 6324
rect 7447 6272 7453 6324
rect 7505 6272 7511 6324
rect 7272 6038 7306 6272
rect 8172 6038 8206 6888
rect 8290 6786 8324 7004
rect 8275 6734 8281 6786
rect 8333 6734 8339 6786
rect 8566 6709 8600 7004
rect 8551 6657 8557 6709
rect 8609 6657 8615 6709
rect 8842 6632 8876 7004
rect 8980 6811 8986 6863
rect 9038 6811 9044 6863
rect 8827 6580 8833 6632
rect 8885 6580 8891 6632
rect 8995 6190 9029 6811
rect 9118 6555 9152 7004
rect 9103 6503 9109 6555
rect 9161 6503 9167 6555
rect 9394 6478 9428 7004
rect 9379 6426 9385 6478
rect 9437 6426 9443 6478
rect 9670 6401 9704 7004
rect 9655 6349 9661 6401
rect 9713 6349 9719 6401
rect 9946 6324 9980 7004
rect 10467 6988 10567 7188
rect 10366 6888 10567 6988
rect 10034 6734 10040 6786
rect 10092 6734 10098 6786
rect 9931 6272 9937 6324
rect 9989 6272 9995 6324
rect 10049 6190 10083 6734
rect 10366 6595 10466 6888
rect 10312 6405 10321 6595
rect 10511 6405 10520 6595
rect 10617 6195 10717 7188
rect 10857 6657 10863 6709
rect 10915 6657 10921 6709
rect 8995 6156 9106 6190
rect 9072 6038 9106 6156
rect 9972 6156 10083 6190
rect 9972 6038 10006 6156
rect 5457 5986 5463 6038
rect 5515 5986 5521 6038
rect 6357 5986 6363 6038
rect 6415 5986 6421 6038
rect 7257 5986 7263 6038
rect 7315 5986 7321 6038
rect 8157 5986 8163 6038
rect 8215 5986 8221 6038
rect 9057 5986 9063 6038
rect 9115 5986 9121 6038
rect 9957 5986 9963 6038
rect 10015 5986 10021 6038
rect 10564 6005 10573 6195
rect 10763 6005 10772 6195
rect 10872 6038 10906 6657
rect 11757 6580 11763 6632
rect 11815 6580 11821 6632
rect 11772 6038 11806 6580
rect 12657 6503 12663 6555
rect 12715 6503 12721 6555
rect 12672 6038 12706 6503
rect 13557 6426 13563 6478
rect 13615 6426 13621 6478
rect 13572 6038 13606 6426
rect 15392 6405 15401 6595
rect 15591 6405 15600 6595
rect 14457 6349 14463 6401
rect 14515 6349 14521 6401
rect 14472 6038 14506 6349
rect 15357 6272 15363 6324
rect 15415 6272 15421 6324
rect 10857 5986 10863 6038
rect 10915 5986 10921 6038
rect 11757 5986 11763 6038
rect 11815 5986 11821 6038
rect 12657 5986 12663 6038
rect 12715 5986 12721 6038
rect 13557 5986 13563 6038
rect 13615 5986 13621 6038
rect 14457 5986 14463 6038
rect 14515 5986 14521 6038
rect 14748 6005 14757 6195
rect 14947 6005 14956 6195
rect 15372 6038 15406 6272
rect 14823 5826 14883 6005
rect 15357 5986 15363 6038
rect 15415 5986 15421 6038
rect 1056 5755 1338 5815
rect 14570 5766 14883 5826
rect 1056 5382 1116 5755
rect 899 5322 1116 5382
rect 14570 5382 14630 5766
rect 14570 5322 14883 5382
rect 899 3072 959 5322
rect 14823 4895 14883 5322
rect 14823 4835 15067 4895
rect 15007 4518 15067 4835
rect 15471 4432 15531 6405
rect 599 595 659 1516
rect 523 405 532 595
rect 722 405 731 595
rect 899 195 959 1816
rect 826 5 835 195
rect 1025 5 1034 195
rect 9864 -342 9898 434
rect 11206 -260 11240 438
rect 12548 -178 12582 434
rect 13890 -96 13924 434
rect 15007 195 15067 1816
rect 15307 595 15367 1516
rect 15234 405 15243 595
rect 15433 405 15442 595
rect 14932 5 14941 195
rect 15131 5 15140 195
rect 16128 -85 16184 -76
rect 13890 -130 16128 -96
rect 16128 -150 16184 -141
rect 16002 -167 16058 -158
rect 12548 -212 16002 -178
rect 16002 -232 16058 -223
rect 16380 -249 16436 -240
rect 11206 -294 16380 -260
rect 16380 -314 16436 -305
rect 16254 -331 16310 -322
rect 9864 -376 16254 -342
rect 16254 -396 16310 -387
<< via2 >>
rect 499 19785 689 19975
rect 16632 20977 16688 21033
rect 16506 20895 16562 20951
rect 16884 20813 16940 20869
rect 16380 20731 16436 20787
rect 16758 20649 16814 20705
rect 14907 19785 15097 19975
rect 799 19385 989 19575
rect 14608 19385 14798 19575
rect 497 15385 687 15575
rect 799 14985 989 15175
rect 4778 14985 4968 15175
rect 5282 15385 5472 15575
rect 10173 15385 10363 15575
rect 14906 15385 15096 15575
rect 10574 14985 10764 15175
rect 14608 14985 14798 15175
rect 5897 14514 5953 14570
rect 6173 14514 6229 14570
rect 6449 14514 6505 14570
rect 6725 14514 6781 14570
rect 7001 14514 7057 14570
rect 7277 14514 7333 14570
rect 7553 14514 7609 14570
rect 7829 14514 7885 14570
rect 8105 14514 8161 14570
rect 8381 14514 8437 14570
rect 8657 14514 8713 14570
rect 8933 14514 8989 14570
rect 9209 14514 9265 14570
rect 9485 14514 9541 14570
rect 9761 14514 9817 14570
rect 10037 14514 10093 14570
rect 5895 14179 5955 14235
rect 6171 14179 6231 14235
rect 6447 14179 6507 14235
rect 6723 14179 6783 14235
rect 6999 14179 7059 14235
rect 7275 14179 7335 14235
rect 7551 14179 7611 14235
rect 7827 14179 7887 14235
rect 8103 14179 8163 14235
rect 8379 14179 8439 14235
rect 8655 14179 8715 14235
rect 8931 14179 8991 14235
rect 9207 14179 9267 14235
rect 9483 14179 9543 14235
rect 9759 14179 9819 14235
rect 10035 14179 10095 14235
rect 5517 7337 5577 7393
rect 5793 7337 5853 7393
rect 6069 7337 6129 7393
rect 6345 7337 6405 7393
rect 6621 7337 6681 7393
rect 6897 7337 6957 7393
rect 7173 7337 7233 7393
rect 7449 7337 7509 7393
rect 7725 7337 7785 7393
rect 8001 7337 8061 7393
rect 8277 7337 8337 7393
rect 8553 7337 8613 7393
rect 8829 7337 8889 7393
rect 9105 7337 9165 7393
rect 9381 7337 9441 7393
rect 9657 7337 9717 7393
rect 9933 7337 9993 7393
rect 5 6405 195 6595
rect 1213 6005 1403 6195
rect 5519 7004 5575 7060
rect 5795 7004 5851 7060
rect 6071 7004 6127 7060
rect 6347 7004 6403 7060
rect 6623 7004 6679 7060
rect 6899 7004 6955 7060
rect 7175 7004 7231 7060
rect 7451 7004 7507 7060
rect 7727 7004 7783 7060
rect 8003 7004 8059 7060
rect 8279 7004 8335 7060
rect 8555 7004 8611 7060
rect 8831 7004 8887 7060
rect 9107 7004 9163 7060
rect 9383 7004 9439 7060
rect 9659 7004 9715 7060
rect 9935 7004 9991 7060
rect 4998 6405 5188 6595
rect 4795 6005 4985 6195
rect 10321 6405 10511 6595
rect 10573 6005 10763 6195
rect 15401 6405 15591 6595
rect 14757 6005 14947 6195
rect 532 405 722 595
rect 835 5 1025 195
rect 15243 405 15433 595
rect 14941 5 15131 195
rect 16128 -141 16184 -85
rect 16002 -223 16058 -167
rect 16380 -305 16436 -249
rect 16254 -387 16310 -331
<< metal3 >>
rect 0 19975 15596 19980
rect 0 19785 499 19975
rect 689 19785 14907 19975
rect 15097 19785 15596 19975
rect 0 19780 15596 19785
rect 0 19575 15596 19580
rect 0 19385 799 19575
rect 989 19385 14608 19575
rect 14798 19385 15596 19575
rect 0 19380 15596 19385
rect 0 15575 15596 15580
rect 0 15385 497 15575
rect 687 15385 5282 15575
rect 5472 15385 10173 15575
rect 10363 15385 14906 15575
rect 15096 15385 15596 15575
rect 0 15380 15596 15385
rect 0 15175 15596 15180
rect 0 14985 799 15175
rect 989 14985 4778 15175
rect 4968 14985 10574 15175
rect 10764 14985 14608 15175
rect 14798 14985 15596 15175
rect 0 14980 15596 14985
rect 5892 14570 5958 14575
rect 5892 14514 5897 14570
rect 5953 14514 5958 14570
rect 5892 14509 5958 14514
rect 6168 14570 6234 14575
rect 6168 14514 6173 14570
rect 6229 14514 6234 14570
rect 6168 14509 6234 14514
rect 6444 14570 6510 14575
rect 6444 14514 6449 14570
rect 6505 14514 6510 14570
rect 6444 14509 6510 14514
rect 6720 14570 6786 14575
rect 6720 14514 6725 14570
rect 6781 14514 6786 14570
rect 6720 14509 6786 14514
rect 6996 14570 7062 14575
rect 6996 14514 7001 14570
rect 7057 14514 7062 14570
rect 6996 14509 7062 14514
rect 7272 14570 7338 14575
rect 7272 14514 7277 14570
rect 7333 14514 7338 14570
rect 7272 14509 7338 14514
rect 7548 14570 7614 14575
rect 7548 14514 7553 14570
rect 7609 14514 7614 14570
rect 7548 14509 7614 14514
rect 7824 14570 7890 14575
rect 7824 14514 7829 14570
rect 7885 14514 7890 14570
rect 7824 14509 7890 14514
rect 8100 14570 8166 14575
rect 8100 14514 8105 14570
rect 8161 14514 8166 14570
rect 8100 14509 8166 14514
rect 8376 14570 8442 14575
rect 8376 14514 8381 14570
rect 8437 14514 8442 14570
rect 8376 14509 8442 14514
rect 8652 14570 8718 14575
rect 8652 14514 8657 14570
rect 8713 14514 8718 14570
rect 8652 14509 8718 14514
rect 8928 14570 8994 14575
rect 8928 14514 8933 14570
rect 8989 14514 8994 14570
rect 8928 14509 8994 14514
rect 9204 14570 9270 14575
rect 9204 14514 9209 14570
rect 9265 14514 9270 14570
rect 9204 14509 9270 14514
rect 9480 14570 9546 14575
rect 9480 14514 9485 14570
rect 9541 14514 9546 14570
rect 9480 14509 9546 14514
rect 9756 14570 9822 14575
rect 9756 14514 9761 14570
rect 9817 14514 9822 14570
rect 9756 14509 9822 14514
rect 10032 14570 10098 14575
rect 10032 14514 10037 14570
rect 10093 14514 10098 14570
rect 10032 14509 10098 14514
rect 5895 14240 5955 14509
rect 6171 14240 6231 14509
rect 6447 14240 6507 14509
rect 6723 14240 6783 14509
rect 6999 14240 7059 14509
rect 7275 14240 7335 14509
rect 7551 14240 7611 14509
rect 7827 14240 7887 14509
rect 8103 14240 8163 14509
rect 8379 14240 8439 14509
rect 8655 14240 8715 14509
rect 8931 14240 8991 14509
rect 9207 14240 9267 14509
rect 9483 14240 9543 14509
rect 9759 14240 9819 14509
rect 10035 14240 10095 14509
rect 5890 14235 5960 14240
rect 5890 14179 5895 14235
rect 5955 14179 5960 14235
rect 5890 14174 5960 14179
rect 6166 14235 6236 14240
rect 6166 14179 6171 14235
rect 6231 14179 6236 14235
rect 6166 14174 6236 14179
rect 6442 14235 6512 14240
rect 6442 14179 6447 14235
rect 6507 14179 6512 14235
rect 6442 14174 6512 14179
rect 6718 14235 6788 14240
rect 6718 14179 6723 14235
rect 6783 14179 6788 14235
rect 6718 14174 6788 14179
rect 6994 14235 7064 14240
rect 6994 14179 6999 14235
rect 7059 14179 7064 14235
rect 6994 14174 7064 14179
rect 7270 14235 7340 14240
rect 7270 14179 7275 14235
rect 7335 14179 7340 14235
rect 7270 14174 7340 14179
rect 7546 14235 7616 14240
rect 7546 14179 7551 14235
rect 7611 14179 7616 14235
rect 7546 14174 7616 14179
rect 7822 14235 7892 14240
rect 7822 14179 7827 14235
rect 7887 14179 7892 14235
rect 7822 14174 7892 14179
rect 8098 14235 8168 14240
rect 8098 14179 8103 14235
rect 8163 14179 8168 14235
rect 8098 14174 8168 14179
rect 8374 14235 8444 14240
rect 8374 14179 8379 14235
rect 8439 14179 8444 14235
rect 8374 14174 8444 14179
rect 8650 14235 8720 14240
rect 8650 14179 8655 14235
rect 8715 14179 8720 14235
rect 8650 14174 8720 14179
rect 8926 14235 8996 14240
rect 8926 14179 8931 14235
rect 8991 14179 8996 14235
rect 8926 14174 8996 14179
rect 9202 14235 9272 14240
rect 9202 14179 9207 14235
rect 9267 14179 9272 14235
rect 9202 14174 9272 14179
rect 9478 14235 9548 14240
rect 9478 14179 9483 14235
rect 9543 14179 9548 14235
rect 9478 14174 9548 14179
rect 9754 14235 9824 14240
rect 9754 14179 9759 14235
rect 9819 14179 9824 14235
rect 9754 14174 9824 14179
rect 10030 14235 10100 14240
rect 10030 14179 10035 14235
rect 10095 14179 10100 14235
rect 10030 14174 10100 14179
rect 5856 13797 10134 13935
rect 5512 7393 5582 7398
rect 5512 7337 5517 7393
rect 5577 7337 5582 7393
rect 5512 7332 5582 7337
rect 5788 7393 5858 7398
rect 5788 7337 5793 7393
rect 5853 7337 5858 7393
rect 5788 7332 5858 7337
rect 6064 7393 6134 7398
rect 6064 7337 6069 7393
rect 6129 7337 6134 7393
rect 6064 7332 6134 7337
rect 6340 7393 6410 7398
rect 6340 7337 6345 7393
rect 6405 7337 6410 7393
rect 6340 7332 6410 7337
rect 6616 7393 6686 7398
rect 6616 7337 6621 7393
rect 6681 7337 6686 7393
rect 6616 7332 6686 7337
rect 6892 7393 6962 7398
rect 6892 7337 6897 7393
rect 6957 7337 6962 7393
rect 6892 7332 6962 7337
rect 7168 7393 7238 7398
rect 7168 7337 7173 7393
rect 7233 7337 7238 7393
rect 7168 7332 7238 7337
rect 7444 7393 7514 7398
rect 7444 7337 7449 7393
rect 7509 7337 7514 7393
rect 7444 7332 7514 7337
rect 7720 7393 7790 7398
rect 7720 7337 7725 7393
rect 7785 7337 7790 7393
rect 7720 7332 7790 7337
rect 7996 7393 8066 7398
rect 7996 7337 8001 7393
rect 8061 7337 8066 7393
rect 7996 7332 8066 7337
rect 8272 7393 8342 7398
rect 8272 7337 8277 7393
rect 8337 7337 8342 7393
rect 8272 7332 8342 7337
rect 8548 7393 8618 7398
rect 8548 7337 8553 7393
rect 8613 7337 8618 7393
rect 8548 7332 8618 7337
rect 8824 7393 8894 7398
rect 8824 7337 8829 7393
rect 8889 7337 8894 7393
rect 8824 7332 8894 7337
rect 9100 7393 9170 7398
rect 9100 7337 9105 7393
rect 9165 7337 9170 7393
rect 9100 7332 9170 7337
rect 9376 7393 9446 7398
rect 9376 7337 9381 7393
rect 9441 7337 9446 7393
rect 9376 7332 9446 7337
rect 9652 7393 9722 7398
rect 9652 7337 9657 7393
rect 9717 7337 9722 7393
rect 9652 7332 9722 7337
rect 9928 7393 9998 7398
rect 9928 7337 9933 7393
rect 9993 7337 9998 7393
rect 9928 7332 9998 7337
rect 5517 7065 5577 7332
rect 5793 7065 5853 7332
rect 6069 7065 6129 7332
rect 6345 7065 6405 7332
rect 6621 7065 6681 7332
rect 6897 7065 6957 7332
rect 7173 7065 7233 7332
rect 7449 7065 7509 7332
rect 7725 7065 7785 7332
rect 8001 7065 8061 7332
rect 8277 7065 8337 7332
rect 8553 7065 8613 7332
rect 8829 7065 8889 7332
rect 9105 7065 9165 7332
rect 9381 7065 9441 7332
rect 9657 7065 9717 7332
rect 9933 7065 9993 7332
rect 5514 7060 5580 7065
rect 5514 7004 5519 7060
rect 5575 7004 5580 7060
rect 5514 6999 5580 7004
rect 5790 7060 5856 7065
rect 5790 7004 5795 7060
rect 5851 7004 5856 7060
rect 5790 6999 5856 7004
rect 6066 7060 6132 7065
rect 6066 7004 6071 7060
rect 6127 7004 6132 7060
rect 6066 6999 6132 7004
rect 6342 7060 6408 7065
rect 6342 7004 6347 7060
rect 6403 7004 6408 7060
rect 6342 6999 6408 7004
rect 6618 7060 6684 7065
rect 6618 7004 6623 7060
rect 6679 7004 6684 7060
rect 6618 6999 6684 7004
rect 6894 7060 6960 7065
rect 6894 7004 6899 7060
rect 6955 7004 6960 7060
rect 6894 6999 6960 7004
rect 7170 7060 7236 7065
rect 7170 7004 7175 7060
rect 7231 7004 7236 7060
rect 7170 6999 7236 7004
rect 7446 7060 7512 7065
rect 7446 7004 7451 7060
rect 7507 7004 7512 7060
rect 7446 6999 7512 7004
rect 7722 7060 7788 7065
rect 7722 7004 7727 7060
rect 7783 7004 7788 7060
rect 7722 6999 7788 7004
rect 7998 7060 8064 7065
rect 7998 7004 8003 7060
rect 8059 7004 8064 7060
rect 7998 6999 8064 7004
rect 8274 7060 8340 7065
rect 8274 7004 8279 7060
rect 8335 7004 8340 7060
rect 8274 6999 8340 7004
rect 8550 7060 8616 7065
rect 8550 7004 8555 7060
rect 8611 7004 8616 7060
rect 8550 6999 8616 7004
rect 8826 7060 8892 7065
rect 8826 7004 8831 7060
rect 8887 7004 8892 7060
rect 8826 6999 8892 7004
rect 9102 7060 9168 7065
rect 9102 7004 9107 7060
rect 9163 7004 9168 7060
rect 9102 6999 9168 7004
rect 9378 7060 9444 7065
rect 9378 7004 9383 7060
rect 9439 7004 9444 7060
rect 9378 6999 9444 7004
rect 9654 7060 9720 7065
rect 9654 7004 9659 7060
rect 9715 7004 9720 7060
rect 9654 6999 9720 7004
rect 9930 7060 9996 7065
rect 9930 7004 9935 7060
rect 9991 7004 9996 7060
rect 9930 6999 9996 7004
rect 0 6595 15596 6600
rect 0 6405 5 6595
rect 195 6405 4998 6595
rect 5188 6405 10321 6595
rect 10511 6405 15401 6595
rect 15591 6405 15596 6595
rect 0 6400 15596 6405
rect 0 6195 15596 6200
rect 0 6005 1213 6195
rect 1403 6005 4795 6195
rect 4985 6005 10573 6195
rect 10763 6005 14757 6195
rect 14947 6005 15596 6195
rect 0 6000 15596 6005
rect 0 595 15596 600
rect 0 405 532 595
rect 722 405 15243 595
rect 15433 405 15596 595
rect 0 400 15596 405
rect 0 195 15596 200
rect 0 5 835 195
rect 1025 5 14941 195
rect 15131 5 15596 195
rect 0 0 15596 5
rect 16000 -162 16060 21433
rect 16126 -80 16186 21433
rect 16123 -85 16189 -80
rect 16123 -141 16128 -85
rect 16184 -141 16189 -85
rect 16123 -146 16189 -141
rect 15997 -167 16063 -162
rect 15997 -223 16002 -167
rect 16058 -223 16063 -167
rect 15997 -228 16063 -223
rect 16252 -326 16312 21433
rect 16378 20792 16438 21433
rect 16504 20956 16564 21433
rect 16630 21038 16690 21433
rect 16627 21033 16693 21038
rect 16627 20977 16632 21033
rect 16688 20977 16693 21033
rect 16627 20972 16693 20977
rect 16501 20951 16567 20956
rect 16501 20895 16506 20951
rect 16562 20895 16567 20951
rect 16501 20890 16567 20895
rect 16375 20787 16441 20792
rect 16375 20731 16380 20787
rect 16436 20731 16441 20787
rect 16375 20726 16441 20731
rect 16378 -244 16438 20726
rect 16504 0 16564 20890
rect 16756 20710 16816 21433
rect 16882 20874 16942 21433
rect 16879 20869 16945 20874
rect 16879 20813 16884 20869
rect 16940 20813 16945 20869
rect 16879 20808 16945 20813
rect 16753 20705 16819 20710
rect 16753 20649 16758 20705
rect 16814 20649 16819 20705
rect 16753 20644 16819 20649
rect 16375 -249 16441 -244
rect 16375 -305 16380 -249
rect 16436 -305 16441 -249
rect 16375 -310 16441 -305
rect 16249 -331 16315 -326
rect 16249 -387 16254 -331
rect 16310 -387 16315 -331
rect 16249 -392 16315 -387
use dac_main  dac_main_0
timestamp 1748333780
transform 1 0 4895 0 1 7088
box 0 0 5822 7394
use lsb_decoder  lsb_decoder_0
timestamp 1748318706
transform 1 0 1128 0 1 15868
box -571 0 13911 4692
use msb_decoder  msb_decoder_0
timestamp 1748318706
transform 1 0 0 0 1 400
box 0 0 15596 5868
<< labels >>
flabel metal3 0 0 15596 200 0 FreeSans 256 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 0 400 15596 600 0 FreeSans 256 0 0 0 VDD
port 2 nsew power bidirectional
flabel metal3 5856 13797 10134 13935 0 FreeSans 256 0 0 0 VOUT
port 3 nsew signal bidirectional
flabel metal3 16882 21133 16942 21433 0 FreeSans 256 0 0 0 IN[0]
port 4 nsew signal input
flabel metal3 16756 21133 16816 21433 0 FreeSans 256 0 0 0 IN[1]
port 5 nsew signal input
flabel metal3 16630 21133 16690 21433 0 FreeSans 256 0 0 0 IN[2]
port 6 nsew signal input
flabel metal3 16504 21133 16564 21433 0 FreeSans 256 0 0 0 IN[3]
port 7 nsew signal input
flabel metal3 16378 21133 16438 21433 0 FreeSans 256 0 0 0 IN[4]
port 8 nsew signal input
flabel metal3 16252 21133 16312 21433 0 FreeSans 256 0 0 0 IN[5]
port 9 nsew signal input
flabel metal3 16126 21133 16186 21433 0 FreeSans 256 0 0 0 IN[6]
port 10 nsew signal input
flabel metal3 16000 21133 16060 21433 0 FreeSans 256 0 0 0 IN[7]
port 11 nsew signal input
<< end >>
