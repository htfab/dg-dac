magic
tech sky130A
magscale 1 2
timestamp 1748318706
<< metal1 >>
rect 0 1132 900 1190
rect 133 99 167 1100
rect 433 99 467 1100
rect 718 534 724 586
rect 776 534 782 586
rect 824 173 858 1017
rect 0 0 900 58
<< via1 >>
rect 724 534 776 586
<< metal2 >>
rect 724 586 776 592
rect 515 543 724 577
rect 724 528 776 534
use inverter_raw  inverter_raw_0
timestamp 1748299149
transform 1 0 512 0 1 -36
box 88 36 388 1226
use nor2_raw  nor2_raw_0
timestamp 1748299149
transform 1 0 -88 0 1 -36
box 88 36 664 1226
<< labels >>
flabel metal1 133 99 167 1100 1 FreeSans 128 0 0 0 A
port 1 n signal input
flabel metal1 433 99 467 1100 1 FreeSans 128 0 0 0 B
port 2 n signal input
flabel metal1 824 173 858 1017 1 FreeSans 128 0 0 0 OUT
port 3 n signal output
flabel metal1 0 0 900 58 1 FreeSans 128 0 0 0 VSS
port 4 n ground bidirectional
flabel metal1 0 1132 900 1190 1 FreeSans 128 0 0 0 VDD
port 5 n power bidirectional
<< end >>
