magic
tech sky130A
magscale 1 2
timestamp 1748337480
<< metal3 >>
rect 7700 32127 7900 32133
rect 14300 32127 14500 32133
rect 20900 32127 21100 32133
rect 6065 31929 7700 32127
rect 7900 31929 14300 32127
rect 14500 31929 20900 32127
rect 21100 31929 21661 32127
rect 6065 31927 21661 31929
rect 7700 31923 7900 31927
rect 14300 31923 14500 31927
rect 20900 31923 21100 31927
rect 7100 31727 7300 31733
rect 13700 31727 13900 31733
rect 20300 31727 20500 31733
rect 6065 31529 7100 31727
rect 7300 31529 13700 31727
rect 13900 31529 20300 31727
rect 20500 31529 21661 31727
rect 6065 31527 21661 31529
rect 7100 31523 7300 31527
rect 13700 31523 13900 31527
rect 20300 31523 20500 31527
rect 6500 31327 6700 31333
rect 13100 31327 13300 31333
rect 19700 31327 19900 31333
rect 6065 31129 6500 31327
rect 6700 31129 13100 31327
rect 13300 31129 19700 31327
rect 19900 31129 21661 31327
rect 6065 31127 21661 31129
rect 6500 31123 6700 31127
rect 13100 31123 13300 31127
rect 19700 31123 19900 31127
<< via3 >>
rect 7700 31929 7900 32127
rect 14300 31929 14500 32127
rect 20900 31929 21100 32127
rect 7100 31529 7300 31727
rect 13700 31529 13900 31727
rect 20300 31529 20500 31727
rect 6500 31129 6700 31327
rect 13100 31129 13300 31327
rect 19700 31129 19900 31327
<< metal4 >>
rect 3006 45015 3066 45152
rect 3558 45015 3618 45152
rect 4110 45015 4170 45152
rect 4662 45015 4722 45152
rect 5214 45015 5274 45152
rect 5766 45015 5826 45152
rect 6318 45015 6378 45152
rect 6870 45015 6930 45152
rect 7422 45015 7482 45152
rect 7974 45015 8034 45152
rect 8526 45015 8586 45152
rect 9078 45015 9138 45152
rect 9630 45015 9690 45152
rect 10182 45015 10242 45152
rect 10734 45015 10794 45152
rect 11286 45015 11346 45152
rect 11838 45015 11898 45152
rect 12390 45015 12450 45152
rect 12942 45015 13002 45152
rect 13494 45015 13554 45152
rect 14046 45015 14106 45152
rect 14598 45015 14658 45152
rect 15150 45015 15210 45152
rect 15702 45015 15762 45152
rect 3003 44949 3069 45015
rect 3555 44949 3621 45015
rect 4107 44949 4173 45015
rect 4659 44949 4725 45015
rect 5211 44949 5277 45015
rect 5763 44949 5829 45015
rect 6315 44949 6381 45015
rect 6867 44949 6933 45015
rect 7419 44949 7485 45015
rect 7971 44949 8037 45015
rect 8523 44949 8589 45015
rect 9075 44949 9141 45015
rect 9627 44949 9693 45015
rect 10179 44949 10245 45015
rect 10731 44949 10797 45015
rect 11283 44949 11349 45015
rect 11835 44949 11901 45015
rect 12387 44949 12453 45015
rect 12939 44949 13005 45015
rect 13491 44949 13557 45015
rect 14043 44949 14109 45015
rect 14595 44949 14661 45015
rect 15147 44949 15213 45015
rect 15699 44949 15765 45015
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 45015 20730 45152
rect 21222 45015 21282 45152
rect 21774 45015 21834 45152
rect 22326 45015 22386 45152
rect 22878 45015 22938 45152
rect 23430 45015 23490 45152
rect 23982 45017 24042 45152
rect 20667 44949 20733 45015
rect 21219 44949 21285 45015
rect 21771 44949 21837 45015
rect 22323 44949 22389 45015
rect 22875 44949 22941 45015
rect 23427 44949 23493 45015
rect 23979 44951 24045 45017
rect 24534 45015 24594 45152
rect 24531 44949 24597 45015
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 6400 31327 6800 44152
rect 6400 31129 6500 31327
rect 6700 31129 6800 31327
rect 6400 1000 6800 31129
rect 7000 31727 7400 44152
rect 7000 31529 7100 31727
rect 7300 31529 7400 31727
rect 7000 1000 7400 31529
rect 7600 32127 8000 44152
rect 7600 31929 7700 32127
rect 7900 31929 8000 32127
rect 7600 1000 8000 31929
rect 13000 31327 13400 44152
rect 13000 31129 13100 31327
rect 13300 31129 13400 31327
rect 13000 1000 13400 31129
rect 13600 31727 14000 44152
rect 13600 31529 13700 31727
rect 13900 31529 14000 31727
rect 13600 1000 14000 31529
rect 14200 32127 14600 44152
rect 14200 31929 14300 32127
rect 14500 31929 14600 32127
rect 14200 1000 14600 31929
rect 19600 31327 20000 44152
rect 19600 31129 19700 31327
rect 19900 31129 20000 31327
rect 19600 1000 20000 31129
rect 20200 31727 20600 44152
rect 20200 31529 20300 31727
rect 20500 31529 20600 31727
rect 20200 1000 20600 31529
rect 20800 32127 21200 44152
rect 20800 31929 20900 32127
rect 21100 31929 21200 32127
rect 20800 1000 21200 31929
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use toplevel_dnwell  toplevel_dnwell_0
timestamp 1748337480
transform 1 0 0 0 1 0
box 0 0 29072 45152
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 6400 1000 6800 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 7000 1000 7400 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 7600 1000 8000 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 19600 1000 20000 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 20200 1000 20600 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 20800 1000 21200 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 13000 1000 13400 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 13600 1000 14000 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 14200 1000 14600 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
