magic
tech sky130A
magscale 1 2
timestamp 1748318706
<< metal1 >>
rect 4807 20196 4813 20248
rect 4865 20196 4871 20248
rect 7503 20196 7509 20248
rect 7561 20196 7567 20248
rect 10199 20196 10205 20248
rect 10257 20196 10263 20248
rect 12595 20202 12601 20254
rect 12653 20202 12659 20254
rect 12895 20196 12901 20248
rect 12953 20196 12959 20248
rect 5899 15680 5951 15686
rect 13776 15680 13828 15686
rect 5951 15637 13776 15671
rect 5899 15622 5951 15628
rect 13776 15622 13828 15628
rect 6175 15603 6227 15609
rect 14473 15603 14525 15609
rect 6227 15560 14473 15594
rect 6175 15545 6227 15551
rect 14473 15545 14525 15551
rect 6451 15526 6503 15532
rect 12434 15526 12486 15532
rect 6503 15483 12434 15517
rect 6451 15468 6503 15474
rect 12434 15468 12486 15474
rect 6727 15449 6779 15455
rect 13131 15449 13183 15455
rect 6779 15406 13131 15440
rect 6727 15391 6779 15397
rect 13131 15391 13183 15397
rect 7003 15372 7055 15378
rect 11092 15372 11144 15378
rect 7055 15329 11092 15363
rect 7003 15314 7055 15320
rect 11092 15314 11144 15320
rect 7279 15295 7331 15301
rect 11789 15295 11841 15301
rect 7331 15252 11789 15286
rect 7279 15237 7331 15243
rect 11789 15237 11841 15243
rect 7555 15218 7607 15224
rect 9750 15218 9802 15224
rect 7607 15175 9750 15209
rect 7555 15160 7607 15166
rect 9750 15160 9802 15166
rect 7831 15141 7883 15147
rect 10447 15141 10499 15147
rect 7883 15098 10447 15132
rect 7831 15083 7883 15089
rect 10447 15083 10499 15089
rect 8107 15064 8159 15070
rect 8482 15064 8534 15070
rect 8159 15021 8482 15055
rect 8107 15006 8159 15012
rect 8482 15006 8534 15012
rect 8383 14987 8435 14993
rect 9105 14987 9157 14993
rect 8435 14944 9105 14978
rect 8383 14929 8435 14935
rect 9105 14929 9157 14935
rect 7140 14910 7192 14916
rect 8659 14910 8711 14916
rect 7192 14867 8659 14901
rect 7140 14852 7192 14858
rect 8659 14852 8711 14858
rect 7689 14833 7741 14839
rect 8935 14833 8987 14839
rect 7741 14790 8935 14824
rect 7689 14775 7741 14781
rect 8935 14775 8987 14781
rect 4382 14756 4434 14762
rect 5724 14756 5776 14762
rect 4434 14713 5510 14747
rect 4382 14698 4434 14704
rect 5079 14679 5131 14685
rect 5131 14636 5433 14670
rect 5079 14621 5131 14627
rect 5399 14516 5433 14636
rect 5476 14593 5510 14713
rect 9211 14756 9263 14762
rect 5776 14713 9211 14747
rect 5724 14698 5776 14704
rect 9211 14698 9263 14704
rect 6347 14679 6399 14685
rect 9487 14679 9539 14685
rect 6399 14636 9487 14670
rect 6347 14621 6399 14627
rect 9487 14621 9539 14627
rect 9763 14602 9815 14608
rect 5476 14559 9763 14593
rect 9763 14544 9815 14550
rect 10039 14525 10091 14531
rect 5399 14482 10039 14516
rect 10039 14467 10091 14473
rect 7729 6940 7781 6946
rect 8163 6940 8215 6946
rect 7781 6897 8163 6931
rect 7729 6882 7781 6888
rect 8163 6882 8215 6888
rect 963 6863 1015 6869
rect 5521 6863 5573 6869
rect 1015 6820 5521 6854
rect 963 6805 1015 6811
rect 5521 6805 5573 6811
rect 8005 6863 8057 6869
rect 8986 6863 9038 6869
rect 8057 6820 8986 6854
rect 8005 6805 8057 6811
rect 8986 6805 9038 6811
rect 1863 6786 1915 6792
rect 5797 6786 5849 6792
rect 1915 6743 5797 6777
rect 1863 6728 1915 6734
rect 5797 6728 5849 6734
rect 8281 6786 8333 6792
rect 10040 6786 10092 6792
rect 8333 6743 10040 6777
rect 8281 6728 8333 6734
rect 10040 6728 10092 6734
rect 2763 6709 2815 6715
rect 6073 6709 6125 6715
rect 2815 6666 6073 6700
rect 2763 6651 2815 6657
rect 6073 6651 6125 6657
rect 8557 6709 8609 6715
rect 10863 6709 10915 6715
rect 8609 6666 10863 6700
rect 8557 6651 8609 6657
rect 10863 6651 10915 6657
rect 3663 6632 3715 6638
rect 6349 6632 6401 6638
rect 3715 6589 6349 6623
rect 3663 6574 3715 6580
rect 6349 6574 6401 6580
rect 8833 6632 8885 6638
rect 11763 6632 11815 6638
rect 8885 6589 11763 6623
rect 8833 6574 8885 6580
rect 11763 6574 11815 6580
rect 4563 6555 4615 6561
rect 6625 6555 6677 6561
rect 4615 6512 6625 6546
rect 4563 6497 4615 6503
rect 6625 6497 6677 6503
rect 9109 6555 9161 6561
rect 12663 6555 12715 6561
rect 9161 6512 12663 6546
rect 9109 6497 9161 6503
rect 12663 6497 12715 6503
rect 5463 6478 5515 6484
rect 6901 6478 6953 6484
rect 5515 6435 6901 6469
rect 5463 6420 5515 6426
rect 6901 6420 6953 6426
rect 9385 6478 9437 6484
rect 13563 6478 13615 6484
rect 9437 6435 13563 6469
rect 9385 6420 9437 6426
rect 13563 6420 13615 6426
rect 6363 6401 6415 6407
rect 7177 6401 7229 6407
rect 6415 6358 7177 6392
rect 6363 6343 6415 6349
rect 7177 6343 7229 6349
rect 9661 6401 9713 6407
rect 14463 6401 14515 6407
rect 9713 6358 14463 6392
rect 9661 6343 9713 6349
rect 14463 6343 14515 6349
rect 7263 6324 7315 6330
rect 7453 6324 7505 6330
rect 7315 6281 7453 6315
rect 7263 6266 7315 6272
rect 7453 6266 7505 6272
rect 9937 6324 9989 6330
rect 15363 6324 15415 6330
rect 9989 6281 15363 6315
rect 9937 6266 9989 6272
rect 15363 6266 15415 6272
rect 963 6038 1015 6044
rect 963 5980 1015 5986
rect 1863 6038 1915 6044
rect 1863 5980 1915 5986
rect 2763 6038 2815 6044
rect 2763 5980 2815 5986
rect 3663 6038 3715 6044
rect 3663 5980 3715 5986
rect 4563 6038 4615 6044
rect 4563 5980 4615 5986
rect 5463 6038 5515 6044
rect 5463 5980 5515 5986
rect 6363 6038 6415 6044
rect 6363 5980 6415 5986
rect 7263 6038 7315 6044
rect 7263 5980 7315 5986
rect 8163 6038 8215 6044
rect 8163 5980 8215 5986
rect 9063 6038 9115 6044
rect 9063 5980 9115 5986
rect 9963 6038 10015 6044
rect 9963 5980 10015 5986
rect 10863 6038 10915 6044
rect 10863 5980 10915 5986
rect 11763 6038 11815 6044
rect 11763 5980 11815 5986
rect 12663 6038 12715 6044
rect 12663 5980 12715 5986
rect 13563 6038 13615 6044
rect 13563 5980 13615 5986
rect 14463 6038 14515 6044
rect 14463 5980 14515 5986
rect 15363 6038 15415 6044
rect 15363 5980 15415 5986
<< via1 >>
rect 4813 20196 4865 20248
rect 7509 20196 7561 20248
rect 10205 20196 10257 20248
rect 12601 20202 12653 20254
rect 12901 20196 12953 20248
rect 5899 15628 5951 15680
rect 13776 15628 13828 15680
rect 6175 15551 6227 15603
rect 14473 15551 14525 15603
rect 6451 15474 6503 15526
rect 12434 15474 12486 15526
rect 6727 15397 6779 15449
rect 13131 15397 13183 15449
rect 7003 15320 7055 15372
rect 11092 15320 11144 15372
rect 7279 15243 7331 15295
rect 11789 15243 11841 15295
rect 7555 15166 7607 15218
rect 9750 15166 9802 15218
rect 7831 15089 7883 15141
rect 10447 15089 10499 15141
rect 8107 15012 8159 15064
rect 8482 15012 8534 15064
rect 8383 14935 8435 14987
rect 9105 14935 9157 14987
rect 7140 14858 7192 14910
rect 8659 14858 8711 14910
rect 7689 14781 7741 14833
rect 8935 14781 8987 14833
rect 4382 14704 4434 14756
rect 5079 14627 5131 14679
rect 5724 14704 5776 14756
rect 9211 14704 9263 14756
rect 6347 14627 6399 14679
rect 9487 14627 9539 14679
rect 9763 14550 9815 14602
rect 10039 14473 10091 14525
rect 7729 6888 7781 6940
rect 8163 6888 8215 6940
rect 963 6811 1015 6863
rect 5521 6811 5573 6863
rect 8005 6811 8057 6863
rect 8986 6811 9038 6863
rect 1863 6734 1915 6786
rect 5797 6734 5849 6786
rect 8281 6734 8333 6786
rect 10040 6734 10092 6786
rect 2763 6657 2815 6709
rect 6073 6657 6125 6709
rect 8557 6657 8609 6709
rect 10863 6657 10915 6709
rect 3663 6580 3715 6632
rect 6349 6580 6401 6632
rect 8833 6580 8885 6632
rect 11763 6580 11815 6632
rect 4563 6503 4615 6555
rect 6625 6503 6677 6555
rect 9109 6503 9161 6555
rect 12663 6503 12715 6555
rect 5463 6426 5515 6478
rect 6901 6426 6953 6478
rect 9385 6426 9437 6478
rect 13563 6426 13615 6478
rect 6363 6349 6415 6401
rect 7177 6349 7229 6401
rect 9661 6349 9713 6401
rect 14463 6349 14515 6401
rect 7263 6272 7315 6324
rect 7453 6272 7505 6324
rect 9937 6272 9989 6324
rect 15363 6272 15415 6324
rect 963 5986 1015 6038
rect 1863 5986 1915 6038
rect 2763 5986 2815 6038
rect 3663 5986 3715 6038
rect 4563 5986 4615 6038
rect 5463 5986 5515 6038
rect 6363 5986 6415 6038
rect 7263 5986 7315 6038
rect 8163 5986 8215 6038
rect 9063 5986 9115 6038
rect 9963 5986 10015 6038
rect 10863 5986 10915 6038
rect 11763 5986 11815 6038
rect 12663 5986 12715 6038
rect 13563 5986 13615 6038
rect 14463 5986 14515 6038
rect 15363 5986 15415 6038
<< metal2 >>
rect 16632 20853 16688 20862
rect 4822 20808 16632 20842
rect 490 19605 499 19795
rect 689 19605 698 19795
rect 564 18473 624 19605
rect 864 19395 924 20285
rect 4822 20254 4856 20808
rect 16632 20788 16688 20797
rect 16506 20771 16562 20780
rect 7518 20726 16506 20760
rect 7518 20254 7552 20726
rect 16506 20706 16562 20715
rect 16884 20689 16940 20698
rect 10214 20644 16884 20678
rect 10214 20254 10248 20644
rect 16884 20624 16940 20633
rect 16380 20607 16436 20616
rect 12610 20562 16380 20596
rect 12610 20260 12644 20562
rect 16380 20542 16436 20551
rect 16758 20525 16814 20534
rect 12910 20480 16758 20514
rect 12601 20254 12653 20260
rect 12910 20254 12944 20480
rect 16758 20460 16814 20469
rect 4813 20248 4865 20254
rect 4813 20190 4865 20196
rect 7509 20248 7561 20254
rect 7509 20190 7561 20196
rect 10205 20248 10257 20254
rect 12601 20196 12653 20202
rect 12901 20248 12953 20254
rect 10205 20190 10257 20196
rect 12901 20190 12953 20196
rect 14672 19395 14732 20285
rect 14898 19605 14907 19795
rect 15097 19605 15106 19795
rect 790 19205 799 19395
rect 989 19205 998 19395
rect 14599 19205 14608 19395
rect 14798 19205 14807 19395
rect 864 18173 924 19205
rect 14672 18173 14732 19205
rect 14972 18473 15032 19605
rect 564 15395 624 16617
rect 488 15205 497 15395
rect 687 15205 696 15395
rect 864 14995 924 16917
rect 790 14805 799 14995
rect 989 14805 998 14995
rect 4391 14756 4425 15800
rect 4769 14805 4778 14995
rect 4968 14805 4977 14995
rect 4376 14704 4382 14756
rect 4434 14704 4440 14756
rect 4823 14504 4923 14805
rect 5088 14679 5122 15800
rect 5273 15205 5282 15395
rect 5472 15205 5481 15395
rect 5073 14627 5079 14679
rect 5131 14627 5137 14679
rect 5327 14504 5427 15205
rect 5733 14756 5767 15800
rect 5893 15628 5899 15680
rect 5951 15628 5957 15680
rect 5718 14704 5724 14756
rect 5776 14704 5782 14756
rect 4823 14404 4995 14504
rect 4895 14202 4995 14404
rect 5045 14404 5427 14504
rect 5045 14202 5145 14404
rect 5908 14390 5942 15628
rect 6169 15551 6175 15603
rect 6227 15551 6233 15603
rect 6430 15594 6464 15800
rect 6356 15560 6464 15594
rect 6184 14390 6218 15551
rect 6356 14679 6390 15560
rect 6445 15474 6451 15526
rect 6503 15474 6509 15526
rect 6341 14627 6347 14679
rect 6399 14627 6405 14679
rect 6460 14390 6494 15474
rect 6721 15397 6727 15449
rect 6779 15397 6785 15449
rect 7075 15440 7109 15800
rect 7075 15406 7183 15440
rect 6736 14390 6770 15397
rect 6997 15320 7003 15372
rect 7055 15320 7061 15372
rect 7012 14390 7046 15320
rect 7149 14910 7183 15406
rect 7273 15243 7279 15295
rect 7331 15243 7337 15295
rect 7134 14858 7140 14910
rect 7192 14858 7198 14910
rect 7288 14390 7322 15243
rect 7549 15166 7555 15218
rect 7607 15166 7613 15218
rect 7772 15209 7806 15800
rect 7698 15175 7806 15209
rect 7564 14390 7598 15166
rect 7698 14833 7732 15175
rect 7825 15089 7831 15141
rect 7883 15089 7889 15141
rect 8417 15132 8451 15800
rect 8417 15098 8525 15132
rect 7683 14781 7689 14833
rect 7741 14781 7747 14833
rect 7840 14390 7874 15089
rect 8491 15064 8525 15098
rect 8101 15012 8107 15064
rect 8159 15012 8165 15064
rect 8476 15012 8482 15064
rect 8534 15012 8540 15064
rect 8116 14390 8150 15012
rect 9114 14987 9148 15800
rect 9759 15218 9793 15800
rect 9744 15166 9750 15218
rect 9802 15166 9808 15218
rect 10164 15205 10173 15395
rect 10363 15205 10372 15395
rect 8377 14935 8383 14987
rect 8435 14935 8441 14987
rect 9099 14935 9105 14987
rect 9157 14935 9163 14987
rect 8392 14390 8426 14935
rect 8653 14858 8659 14910
rect 8711 14858 8717 14910
rect 8668 14390 8702 14858
rect 8929 14781 8935 14833
rect 8987 14781 8993 14833
rect 8944 14390 8978 14781
rect 9205 14704 9211 14756
rect 9263 14704 9269 14756
rect 10218 14704 10318 15205
rect 10456 15141 10490 15800
rect 11101 15372 11135 15800
rect 11086 15320 11092 15372
rect 11144 15320 11150 15372
rect 11798 15295 11832 15800
rect 12443 15526 12477 15800
rect 12428 15474 12434 15526
rect 12486 15474 12492 15526
rect 13140 15449 13174 15800
rect 13785 15680 13819 15800
rect 13770 15628 13776 15680
rect 13828 15628 13834 15680
rect 14482 15603 14516 15800
rect 14467 15551 14473 15603
rect 14525 15551 14531 15603
rect 13125 15397 13131 15449
rect 13183 15397 13189 15449
rect 11783 15243 11789 15295
rect 11841 15243 11847 15295
rect 10441 15089 10447 15141
rect 10499 15089 10505 15141
rect 14672 14995 14732 16917
rect 14972 15395 15032 16617
rect 14897 15205 14906 15395
rect 15096 15205 15105 15395
rect 10565 14805 10574 14995
rect 10764 14805 10773 14995
rect 14599 14805 14608 14995
rect 14798 14805 14807 14995
rect 9220 14390 9254 14704
rect 9481 14627 9487 14679
rect 9539 14627 9545 14679
rect 9496 14390 9530 14627
rect 10218 14604 10567 14704
rect 9757 14550 9763 14602
rect 9815 14550 9821 14602
rect 9772 14390 9806 14550
rect 10033 14473 10039 14525
rect 10091 14473 10097 14525
rect 10048 14390 10082 14473
rect 5888 14334 5897 14390
rect 5953 14334 5962 14390
rect 6164 14334 6173 14390
rect 6229 14334 6238 14390
rect 6440 14334 6449 14390
rect 6505 14334 6514 14390
rect 6716 14334 6725 14390
rect 6781 14334 6790 14390
rect 6992 14334 7001 14390
rect 7057 14334 7066 14390
rect 7268 14334 7277 14390
rect 7333 14334 7342 14390
rect 7544 14334 7553 14390
rect 7609 14334 7618 14390
rect 7820 14334 7829 14390
rect 7885 14334 7894 14390
rect 8096 14334 8105 14390
rect 8161 14334 8170 14390
rect 8372 14334 8381 14390
rect 8437 14334 8446 14390
rect 8648 14334 8657 14390
rect 8713 14334 8722 14390
rect 8924 14334 8933 14390
rect 8989 14334 8998 14390
rect 9200 14334 9209 14390
rect 9265 14334 9274 14390
rect 9476 14334 9485 14390
rect 9541 14334 9550 14390
rect 9752 14334 9761 14390
rect 9817 14334 9826 14390
rect 10028 14334 10037 14390
rect 10093 14334 10102 14390
rect 10467 14202 10567 14604
rect 10617 14202 10717 14805
rect 5895 14055 5955 14064
rect 5895 13828 5955 13999
rect 6171 14055 6231 14064
rect 6171 13828 6231 13999
rect 6447 14055 6507 14064
rect 6447 13828 6507 13999
rect 6723 14055 6783 14064
rect 6723 13828 6783 13999
rect 6999 14055 7059 14064
rect 6999 13828 7059 13999
rect 7275 14055 7335 14064
rect 7275 13828 7335 13999
rect 7551 14055 7611 14064
rect 7551 13828 7611 13999
rect 7827 14055 7887 14064
rect 7827 13828 7887 13999
rect 8103 14055 8163 14064
rect 8103 13828 8163 13999
rect 8379 14055 8439 14064
rect 8379 13828 8439 13999
rect 8655 14055 8715 14064
rect 8655 13828 8715 13999
rect 8931 14055 8991 14064
rect 8931 13828 8991 13999
rect 9207 14055 9267 14064
rect 9207 13828 9267 13999
rect 9483 14055 9543 14064
rect 9483 13828 9543 13999
rect 9759 14055 9819 14064
rect 9759 13828 9819 13999
rect 10035 14055 10095 14064
rect 10035 13828 10095 13999
rect 5517 7393 5577 7562
rect 5517 7328 5577 7337
rect 5793 7393 5853 7562
rect 5793 7328 5853 7337
rect 6069 7393 6129 7562
rect 6069 7328 6129 7337
rect 6345 7393 6405 7562
rect 6345 7328 6405 7337
rect 6621 7393 6681 7562
rect 6621 7328 6681 7337
rect 6897 7393 6957 7562
rect 6897 7328 6957 7337
rect 7173 7393 7233 7562
rect 7173 7328 7233 7337
rect 7449 7393 7509 7562
rect 7449 7328 7509 7337
rect 7725 7393 7785 7562
rect 7725 7328 7785 7337
rect 8001 7393 8061 7562
rect 8001 7328 8061 7337
rect 8277 7393 8337 7562
rect 8277 7328 8337 7337
rect 8553 7393 8613 7562
rect 8553 7328 8613 7337
rect 8829 7393 8889 7562
rect 8829 7328 8889 7337
rect 9105 7393 9165 7562
rect 9105 7328 9165 7337
rect 9381 7393 9441 7562
rect 9381 7328 9441 7337
rect 9657 7393 9717 7562
rect 9657 7328 9717 7337
rect 9933 7393 9993 7562
rect 9933 7328 9993 7337
rect 4840 7088 4995 7188
rect 957 6811 963 6863
rect 1015 6811 1021 6863
rect -4 6405 5 6595
rect 195 6405 204 6595
rect 65 4432 125 6405
rect 972 6038 1006 6811
rect 1857 6734 1863 6786
rect 1915 6734 1921 6786
rect 957 5986 963 6038
rect 1015 5986 1021 6038
rect 1204 6005 1213 6195
rect 1403 6005 1412 6195
rect 1872 6038 1906 6734
rect 2757 6657 2763 6709
rect 2815 6657 2821 6709
rect 2772 6038 2806 6657
rect 3657 6580 3663 6632
rect 3715 6580 3721 6632
rect 3672 6038 3706 6580
rect 4557 6503 4563 6555
rect 4615 6503 4621 6555
rect 4572 6038 4606 6503
rect 4840 6195 4940 7088
rect 5045 6595 5145 7188
rect 5510 7004 5519 7060
rect 5575 7004 5584 7060
rect 5786 7004 5795 7060
rect 5851 7004 5860 7060
rect 6062 7004 6071 7060
rect 6127 7004 6136 7060
rect 6338 7004 6347 7060
rect 6403 7004 6412 7060
rect 6614 7004 6623 7060
rect 6679 7004 6688 7060
rect 6890 7004 6899 7060
rect 6955 7004 6964 7060
rect 7166 7004 7175 7060
rect 7231 7004 7240 7060
rect 7442 7004 7451 7060
rect 7507 7004 7516 7060
rect 7718 7004 7727 7060
rect 7783 7004 7792 7060
rect 7994 7004 8003 7060
rect 8059 7004 8068 7060
rect 8270 7004 8279 7060
rect 8335 7004 8344 7060
rect 8546 7004 8555 7060
rect 8611 7004 8620 7060
rect 8822 7004 8831 7060
rect 8887 7004 8896 7060
rect 9098 7004 9107 7060
rect 9163 7004 9172 7060
rect 9374 7004 9383 7060
rect 9439 7004 9448 7060
rect 9650 7004 9659 7060
rect 9715 7004 9724 7060
rect 9926 7004 9935 7060
rect 9991 7004 10000 7060
rect 5530 6863 5564 7004
rect 5515 6811 5521 6863
rect 5573 6811 5579 6863
rect 5806 6786 5840 7004
rect 5791 6734 5797 6786
rect 5849 6734 5855 6786
rect 6082 6709 6116 7004
rect 6067 6657 6073 6709
rect 6125 6657 6131 6709
rect 6358 6632 6392 7004
rect 4989 6405 4998 6595
rect 5188 6405 5197 6595
rect 6343 6580 6349 6632
rect 6401 6580 6407 6632
rect 6634 6555 6668 7004
rect 6619 6503 6625 6555
rect 6677 6503 6683 6555
rect 6910 6478 6944 7004
rect 5457 6426 5463 6478
rect 5515 6426 5521 6478
rect 6895 6426 6901 6478
rect 6953 6426 6959 6478
rect 1278 5815 1338 6005
rect 1857 5986 1863 6038
rect 1915 5986 1921 6038
rect 2757 5986 2763 6038
rect 2815 5986 2821 6038
rect 3657 5986 3663 6038
rect 3715 5986 3721 6038
rect 4557 5986 4563 6038
rect 4615 5986 4621 6038
rect 4786 6005 4795 6195
rect 4985 6005 4994 6195
rect 5472 6038 5506 6426
rect 7186 6401 7220 7004
rect 6357 6349 6363 6401
rect 6415 6349 6421 6401
rect 7171 6349 7177 6401
rect 7229 6349 7235 6401
rect 6372 6038 6406 6349
rect 7462 6324 7496 7004
rect 7738 6940 7772 7004
rect 7723 6888 7729 6940
rect 7781 6888 7787 6940
rect 8014 6863 8048 7004
rect 8157 6888 8163 6940
rect 8215 6888 8221 6940
rect 7999 6811 8005 6863
rect 8057 6811 8063 6863
rect 7257 6272 7263 6324
rect 7315 6272 7321 6324
rect 7447 6272 7453 6324
rect 7505 6272 7511 6324
rect 7272 6038 7306 6272
rect 8172 6038 8206 6888
rect 8290 6786 8324 7004
rect 8275 6734 8281 6786
rect 8333 6734 8339 6786
rect 8566 6709 8600 7004
rect 8551 6657 8557 6709
rect 8609 6657 8615 6709
rect 8842 6632 8876 7004
rect 8980 6811 8986 6863
rect 9038 6811 9044 6863
rect 8827 6580 8833 6632
rect 8885 6580 8891 6632
rect 8995 6190 9029 6811
rect 9118 6555 9152 7004
rect 9103 6503 9109 6555
rect 9161 6503 9167 6555
rect 9394 6478 9428 7004
rect 9379 6426 9385 6478
rect 9437 6426 9443 6478
rect 9670 6401 9704 7004
rect 9655 6349 9661 6401
rect 9713 6349 9719 6401
rect 9946 6324 9980 7004
rect 10467 6988 10567 7188
rect 10366 6888 10567 6988
rect 10034 6734 10040 6786
rect 10092 6734 10098 6786
rect 9931 6272 9937 6324
rect 9989 6272 9995 6324
rect 10049 6190 10083 6734
rect 10366 6595 10466 6888
rect 10312 6405 10321 6595
rect 10511 6405 10520 6595
rect 10617 6195 10717 7188
rect 10857 6657 10863 6709
rect 10915 6657 10921 6709
rect 8995 6156 9106 6190
rect 9072 6038 9106 6156
rect 9972 6156 10083 6190
rect 9972 6038 10006 6156
rect 5457 5986 5463 6038
rect 5515 5986 5521 6038
rect 6357 5986 6363 6038
rect 6415 5986 6421 6038
rect 7257 5986 7263 6038
rect 7315 5986 7321 6038
rect 8157 5986 8163 6038
rect 8215 5986 8221 6038
rect 9057 5986 9063 6038
rect 9115 5986 9121 6038
rect 9957 5986 9963 6038
rect 10015 5986 10021 6038
rect 10564 6005 10573 6195
rect 10763 6005 10772 6195
rect 10872 6038 10906 6657
rect 11757 6580 11763 6632
rect 11815 6580 11821 6632
rect 11772 6038 11806 6580
rect 12657 6503 12663 6555
rect 12715 6503 12721 6555
rect 12672 6038 12706 6503
rect 13557 6426 13563 6478
rect 13615 6426 13621 6478
rect 13572 6038 13606 6426
rect 15392 6405 15401 6595
rect 15591 6405 15600 6595
rect 14457 6349 14463 6401
rect 14515 6349 14521 6401
rect 14472 6038 14506 6349
rect 15357 6272 15363 6324
rect 15415 6272 15421 6324
rect 10857 5986 10863 6038
rect 10915 5986 10921 6038
rect 11757 5986 11763 6038
rect 11815 5986 11821 6038
rect 12657 5986 12663 6038
rect 12715 5986 12721 6038
rect 13557 5986 13563 6038
rect 13615 5986 13621 6038
rect 14457 5986 14463 6038
rect 14515 5986 14521 6038
rect 14748 6005 14757 6195
rect 14947 6005 14956 6195
rect 15372 6038 15406 6272
rect 14823 5826 14883 6005
rect 15357 5986 15363 6038
rect 15415 5986 15421 6038
rect 1056 5755 1338 5815
rect 14570 5766 14883 5826
rect 1056 5382 1116 5755
rect 899 5322 1116 5382
rect 14570 5382 14630 5766
rect 14570 5322 14883 5382
rect 899 3072 959 5322
rect 14823 4895 14883 5322
rect 14823 4835 15067 4895
rect 15007 4518 15067 4835
rect 15471 4432 15531 6405
rect 599 595 659 1516
rect 523 405 532 595
rect 722 405 731 595
rect 899 195 959 1816
rect 826 5 835 195
rect 1025 5 1034 195
rect 9864 -342 9898 434
rect 11206 -260 11240 438
rect 12548 -178 12582 434
rect 13890 -96 13924 434
rect 15007 195 15067 1816
rect 15307 595 15367 1516
rect 15234 405 15243 595
rect 15433 405 15442 595
rect 14932 5 14941 195
rect 15131 5 15140 195
rect 16128 -85 16184 -76
rect 13890 -130 16128 -96
rect 16128 -150 16184 -141
rect 16002 -167 16058 -158
rect 12548 -212 16002 -178
rect 16002 -232 16058 -223
rect 16380 -249 16436 -240
rect 11206 -294 16380 -260
rect 16380 -314 16436 -305
rect 16254 -331 16310 -322
rect 9864 -376 16254 -342
rect 16254 -396 16310 -387
<< via2 >>
rect 499 19605 689 19795
rect 16632 20797 16688 20853
rect 16506 20715 16562 20771
rect 16884 20633 16940 20689
rect 16380 20551 16436 20607
rect 16758 20469 16814 20525
rect 14907 19605 15097 19795
rect 799 19205 989 19395
rect 14608 19205 14798 19395
rect 497 15205 687 15395
rect 799 14805 989 14995
rect 4778 14805 4968 14995
rect 5282 15205 5472 15395
rect 10173 15205 10363 15395
rect 14906 15205 15096 15395
rect 10574 14805 10764 14995
rect 14608 14805 14798 14995
rect 5897 14334 5953 14390
rect 6173 14334 6229 14390
rect 6449 14334 6505 14390
rect 6725 14334 6781 14390
rect 7001 14334 7057 14390
rect 7277 14334 7333 14390
rect 7553 14334 7609 14390
rect 7829 14334 7885 14390
rect 8105 14334 8161 14390
rect 8381 14334 8437 14390
rect 8657 14334 8713 14390
rect 8933 14334 8989 14390
rect 9209 14334 9265 14390
rect 9485 14334 9541 14390
rect 9761 14334 9817 14390
rect 10037 14334 10093 14390
rect 5895 13999 5955 14055
rect 6171 13999 6231 14055
rect 6447 13999 6507 14055
rect 6723 13999 6783 14055
rect 6999 13999 7059 14055
rect 7275 13999 7335 14055
rect 7551 13999 7611 14055
rect 7827 13999 7887 14055
rect 8103 13999 8163 14055
rect 8379 13999 8439 14055
rect 8655 13999 8715 14055
rect 8931 13999 8991 14055
rect 9207 13999 9267 14055
rect 9483 13999 9543 14055
rect 9759 13999 9819 14055
rect 10035 13999 10095 14055
rect 5517 7337 5577 7393
rect 5793 7337 5853 7393
rect 6069 7337 6129 7393
rect 6345 7337 6405 7393
rect 6621 7337 6681 7393
rect 6897 7337 6957 7393
rect 7173 7337 7233 7393
rect 7449 7337 7509 7393
rect 7725 7337 7785 7393
rect 8001 7337 8061 7393
rect 8277 7337 8337 7393
rect 8553 7337 8613 7393
rect 8829 7337 8889 7393
rect 9105 7337 9165 7393
rect 9381 7337 9441 7393
rect 9657 7337 9717 7393
rect 9933 7337 9993 7393
rect 5 6405 195 6595
rect 1213 6005 1403 6195
rect 5519 7004 5575 7060
rect 5795 7004 5851 7060
rect 6071 7004 6127 7060
rect 6347 7004 6403 7060
rect 6623 7004 6679 7060
rect 6899 7004 6955 7060
rect 7175 7004 7231 7060
rect 7451 7004 7507 7060
rect 7727 7004 7783 7060
rect 8003 7004 8059 7060
rect 8279 7004 8335 7060
rect 8555 7004 8611 7060
rect 8831 7004 8887 7060
rect 9107 7004 9163 7060
rect 9383 7004 9439 7060
rect 9659 7004 9715 7060
rect 9935 7004 9991 7060
rect 4998 6405 5188 6595
rect 4795 6005 4985 6195
rect 10321 6405 10511 6595
rect 10573 6005 10763 6195
rect 15401 6405 15591 6595
rect 14757 6005 14947 6195
rect 532 405 722 595
rect 835 5 1025 195
rect 15243 405 15433 595
rect 14941 5 15131 195
rect 16128 -141 16184 -85
rect 16002 -223 16058 -167
rect 16380 -305 16436 -249
rect 16254 -387 16310 -331
<< metal3 >>
rect 0 19795 15596 19800
rect 0 19605 499 19795
rect 689 19605 14907 19795
rect 15097 19605 15596 19795
rect 0 19600 15596 19605
rect 0 19395 15596 19400
rect 0 19205 799 19395
rect 989 19205 14608 19395
rect 14798 19205 15596 19395
rect 0 19200 15596 19205
rect 0 15395 15596 15400
rect 0 15205 497 15395
rect 687 15205 5282 15395
rect 5472 15205 10173 15395
rect 10363 15205 14906 15395
rect 15096 15205 15596 15395
rect 0 15200 15596 15205
rect 0 14995 15596 15000
rect 0 14805 799 14995
rect 989 14805 4778 14995
rect 4968 14805 10574 14995
rect 10764 14805 14608 14995
rect 14798 14805 15596 14995
rect 0 14800 15596 14805
rect 5892 14390 5958 14395
rect 5892 14334 5897 14390
rect 5953 14334 5958 14390
rect 5892 14329 5958 14334
rect 6168 14390 6234 14395
rect 6168 14334 6173 14390
rect 6229 14334 6234 14390
rect 6168 14329 6234 14334
rect 6444 14390 6510 14395
rect 6444 14334 6449 14390
rect 6505 14334 6510 14390
rect 6444 14329 6510 14334
rect 6720 14390 6786 14395
rect 6720 14334 6725 14390
rect 6781 14334 6786 14390
rect 6720 14329 6786 14334
rect 6996 14390 7062 14395
rect 6996 14334 7001 14390
rect 7057 14334 7062 14390
rect 6996 14329 7062 14334
rect 7272 14390 7338 14395
rect 7272 14334 7277 14390
rect 7333 14334 7338 14390
rect 7272 14329 7338 14334
rect 7548 14390 7614 14395
rect 7548 14334 7553 14390
rect 7609 14334 7614 14390
rect 7548 14329 7614 14334
rect 7824 14390 7890 14395
rect 7824 14334 7829 14390
rect 7885 14334 7890 14390
rect 7824 14329 7890 14334
rect 8100 14390 8166 14395
rect 8100 14334 8105 14390
rect 8161 14334 8166 14390
rect 8100 14329 8166 14334
rect 8376 14390 8442 14395
rect 8376 14334 8381 14390
rect 8437 14334 8442 14390
rect 8376 14329 8442 14334
rect 8652 14390 8718 14395
rect 8652 14334 8657 14390
rect 8713 14334 8718 14390
rect 8652 14329 8718 14334
rect 8928 14390 8994 14395
rect 8928 14334 8933 14390
rect 8989 14334 8994 14390
rect 8928 14329 8994 14334
rect 9204 14390 9270 14395
rect 9204 14334 9209 14390
rect 9265 14334 9270 14390
rect 9204 14329 9270 14334
rect 9480 14390 9546 14395
rect 9480 14334 9485 14390
rect 9541 14334 9546 14390
rect 9480 14329 9546 14334
rect 9756 14390 9822 14395
rect 9756 14334 9761 14390
rect 9817 14334 9822 14390
rect 9756 14329 9822 14334
rect 10032 14390 10098 14395
rect 10032 14334 10037 14390
rect 10093 14334 10098 14390
rect 10032 14329 10098 14334
rect 5895 14060 5955 14329
rect 6171 14060 6231 14329
rect 6447 14060 6507 14329
rect 6723 14060 6783 14329
rect 6999 14060 7059 14329
rect 7275 14060 7335 14329
rect 7551 14060 7611 14329
rect 7827 14060 7887 14329
rect 8103 14060 8163 14329
rect 8379 14060 8439 14329
rect 8655 14060 8715 14329
rect 8931 14060 8991 14329
rect 9207 14060 9267 14329
rect 9483 14060 9543 14329
rect 9759 14060 9819 14329
rect 10035 14060 10095 14329
rect 5890 14055 5960 14060
rect 5890 13999 5895 14055
rect 5955 13999 5960 14055
rect 5890 13994 5960 13999
rect 6166 14055 6236 14060
rect 6166 13999 6171 14055
rect 6231 13999 6236 14055
rect 6166 13994 6236 13999
rect 6442 14055 6512 14060
rect 6442 13999 6447 14055
rect 6507 13999 6512 14055
rect 6442 13994 6512 13999
rect 6718 14055 6788 14060
rect 6718 13999 6723 14055
rect 6783 13999 6788 14055
rect 6718 13994 6788 13999
rect 6994 14055 7064 14060
rect 6994 13999 6999 14055
rect 7059 13999 7064 14055
rect 6994 13994 7064 13999
rect 7270 14055 7340 14060
rect 7270 13999 7275 14055
rect 7335 13999 7340 14055
rect 7270 13994 7340 13999
rect 7546 14055 7616 14060
rect 7546 13999 7551 14055
rect 7611 13999 7616 14055
rect 7546 13994 7616 13999
rect 7822 14055 7892 14060
rect 7822 13999 7827 14055
rect 7887 13999 7892 14055
rect 7822 13994 7892 13999
rect 8098 14055 8168 14060
rect 8098 13999 8103 14055
rect 8163 13999 8168 14055
rect 8098 13994 8168 13999
rect 8374 14055 8444 14060
rect 8374 13999 8379 14055
rect 8439 13999 8444 14055
rect 8374 13994 8444 13999
rect 8650 14055 8720 14060
rect 8650 13999 8655 14055
rect 8715 13999 8720 14055
rect 8650 13994 8720 13999
rect 8926 14055 8996 14060
rect 8926 13999 8931 14055
rect 8991 13999 8996 14055
rect 8926 13994 8996 13999
rect 9202 14055 9272 14060
rect 9202 13999 9207 14055
rect 9267 13999 9272 14055
rect 9202 13994 9272 13999
rect 9478 14055 9548 14060
rect 9478 13999 9483 14055
rect 9543 13999 9548 14055
rect 9478 13994 9548 13999
rect 9754 14055 9824 14060
rect 9754 13999 9759 14055
rect 9819 13999 9824 14055
rect 9754 13994 9824 13999
rect 10030 14055 10100 14060
rect 10030 13999 10035 14055
rect 10095 13999 10100 14055
rect 10030 13994 10100 13999
rect 5856 13617 10134 13755
rect 5512 7393 5582 7398
rect 5512 7337 5517 7393
rect 5577 7337 5582 7393
rect 5512 7332 5582 7337
rect 5788 7393 5858 7398
rect 5788 7337 5793 7393
rect 5853 7337 5858 7393
rect 5788 7332 5858 7337
rect 6064 7393 6134 7398
rect 6064 7337 6069 7393
rect 6129 7337 6134 7393
rect 6064 7332 6134 7337
rect 6340 7393 6410 7398
rect 6340 7337 6345 7393
rect 6405 7337 6410 7393
rect 6340 7332 6410 7337
rect 6616 7393 6686 7398
rect 6616 7337 6621 7393
rect 6681 7337 6686 7393
rect 6616 7332 6686 7337
rect 6892 7393 6962 7398
rect 6892 7337 6897 7393
rect 6957 7337 6962 7393
rect 6892 7332 6962 7337
rect 7168 7393 7238 7398
rect 7168 7337 7173 7393
rect 7233 7337 7238 7393
rect 7168 7332 7238 7337
rect 7444 7393 7514 7398
rect 7444 7337 7449 7393
rect 7509 7337 7514 7393
rect 7444 7332 7514 7337
rect 7720 7393 7790 7398
rect 7720 7337 7725 7393
rect 7785 7337 7790 7393
rect 7720 7332 7790 7337
rect 7996 7393 8066 7398
rect 7996 7337 8001 7393
rect 8061 7337 8066 7393
rect 7996 7332 8066 7337
rect 8272 7393 8342 7398
rect 8272 7337 8277 7393
rect 8337 7337 8342 7393
rect 8272 7332 8342 7337
rect 8548 7393 8618 7398
rect 8548 7337 8553 7393
rect 8613 7337 8618 7393
rect 8548 7332 8618 7337
rect 8824 7393 8894 7398
rect 8824 7337 8829 7393
rect 8889 7337 8894 7393
rect 8824 7332 8894 7337
rect 9100 7393 9170 7398
rect 9100 7337 9105 7393
rect 9165 7337 9170 7393
rect 9100 7332 9170 7337
rect 9376 7393 9446 7398
rect 9376 7337 9381 7393
rect 9441 7337 9446 7393
rect 9376 7332 9446 7337
rect 9652 7393 9722 7398
rect 9652 7337 9657 7393
rect 9717 7337 9722 7393
rect 9652 7332 9722 7337
rect 9928 7393 9998 7398
rect 9928 7337 9933 7393
rect 9993 7337 9998 7393
rect 9928 7332 9998 7337
rect 5517 7065 5577 7332
rect 5793 7065 5853 7332
rect 6069 7065 6129 7332
rect 6345 7065 6405 7332
rect 6621 7065 6681 7332
rect 6897 7065 6957 7332
rect 7173 7065 7233 7332
rect 7449 7065 7509 7332
rect 7725 7065 7785 7332
rect 8001 7065 8061 7332
rect 8277 7065 8337 7332
rect 8553 7065 8613 7332
rect 8829 7065 8889 7332
rect 9105 7065 9165 7332
rect 9381 7065 9441 7332
rect 9657 7065 9717 7332
rect 9933 7065 9993 7332
rect 5514 7060 5580 7065
rect 5514 7004 5519 7060
rect 5575 7004 5580 7060
rect 5514 6999 5580 7004
rect 5790 7060 5856 7065
rect 5790 7004 5795 7060
rect 5851 7004 5856 7060
rect 5790 6999 5856 7004
rect 6066 7060 6132 7065
rect 6066 7004 6071 7060
rect 6127 7004 6132 7060
rect 6066 6999 6132 7004
rect 6342 7060 6408 7065
rect 6342 7004 6347 7060
rect 6403 7004 6408 7060
rect 6342 6999 6408 7004
rect 6618 7060 6684 7065
rect 6618 7004 6623 7060
rect 6679 7004 6684 7060
rect 6618 6999 6684 7004
rect 6894 7060 6960 7065
rect 6894 7004 6899 7060
rect 6955 7004 6960 7060
rect 6894 6999 6960 7004
rect 7170 7060 7236 7065
rect 7170 7004 7175 7060
rect 7231 7004 7236 7060
rect 7170 6999 7236 7004
rect 7446 7060 7512 7065
rect 7446 7004 7451 7060
rect 7507 7004 7512 7060
rect 7446 6999 7512 7004
rect 7722 7060 7788 7065
rect 7722 7004 7727 7060
rect 7783 7004 7788 7060
rect 7722 6999 7788 7004
rect 7998 7060 8064 7065
rect 7998 7004 8003 7060
rect 8059 7004 8064 7060
rect 7998 6999 8064 7004
rect 8274 7060 8340 7065
rect 8274 7004 8279 7060
rect 8335 7004 8340 7060
rect 8274 6999 8340 7004
rect 8550 7060 8616 7065
rect 8550 7004 8555 7060
rect 8611 7004 8616 7060
rect 8550 6999 8616 7004
rect 8826 7060 8892 7065
rect 8826 7004 8831 7060
rect 8887 7004 8892 7060
rect 8826 6999 8892 7004
rect 9102 7060 9168 7065
rect 9102 7004 9107 7060
rect 9163 7004 9168 7060
rect 9102 6999 9168 7004
rect 9378 7060 9444 7065
rect 9378 7004 9383 7060
rect 9439 7004 9444 7060
rect 9378 6999 9444 7004
rect 9654 7060 9720 7065
rect 9654 7004 9659 7060
rect 9715 7004 9720 7060
rect 9654 6999 9720 7004
rect 9930 7060 9996 7065
rect 9930 7004 9935 7060
rect 9991 7004 9996 7060
rect 9930 6999 9996 7004
rect 0 6595 15596 6600
rect 0 6405 5 6595
rect 195 6405 4998 6595
rect 5188 6405 10321 6595
rect 10511 6405 15401 6595
rect 15591 6405 15596 6595
rect 0 6400 15596 6405
rect 0 6195 15596 6200
rect 0 6005 1213 6195
rect 1403 6005 4795 6195
rect 4985 6005 10573 6195
rect 10763 6005 14757 6195
rect 14947 6005 15596 6195
rect 0 6000 15596 6005
rect 0 595 15596 600
rect 0 405 532 595
rect 722 405 15243 595
rect 15433 405 15596 595
rect 0 400 15596 405
rect 0 195 15596 200
rect 0 5 835 195
rect 1025 5 14941 195
rect 15131 5 15596 195
rect 0 0 15596 5
rect 16000 -162 16060 21253
rect 16126 -80 16186 21253
rect 16123 -85 16189 -80
rect 16123 -141 16128 -85
rect 16184 -141 16189 -85
rect 16123 -146 16189 -141
rect 15997 -167 16063 -162
rect 15997 -223 16002 -167
rect 16058 -223 16063 -167
rect 15997 -228 16063 -223
rect 16252 -326 16312 21253
rect 16378 20612 16438 21253
rect 16504 20776 16564 21253
rect 16630 20858 16690 21253
rect 16627 20853 16693 20858
rect 16627 20797 16632 20853
rect 16688 20797 16693 20853
rect 16627 20792 16693 20797
rect 16501 20771 16567 20776
rect 16501 20715 16506 20771
rect 16562 20715 16567 20771
rect 16501 20710 16567 20715
rect 16375 20607 16441 20612
rect 16375 20551 16380 20607
rect 16436 20551 16441 20607
rect 16375 20546 16441 20551
rect 16378 -244 16438 20546
rect 16504 0 16564 20710
rect 16756 20530 16816 21253
rect 16882 20694 16942 21253
rect 16879 20689 16945 20694
rect 16879 20633 16884 20689
rect 16940 20633 16945 20689
rect 16879 20628 16945 20633
rect 16753 20525 16819 20530
rect 16753 20469 16758 20525
rect 16814 20469 16819 20525
rect 16753 20464 16819 20469
rect 16375 -249 16441 -244
rect 16375 -305 16380 -249
rect 16436 -305 16441 -249
rect 16375 -310 16441 -305
rect 16249 -331 16315 -326
rect 16249 -387 16254 -331
rect 16310 -387 16315 -331
rect 16249 -392 16315 -387
use dac_main  dac_main_0
timestamp 1748309517
transform 1 0 4895 0 1 7088
box 0 0 5822 7214
use lsb_decoder  lsb_decoder_0
timestamp 1748318706
transform 1 0 1128 0 1 15688
box -571 0 13911 4692
use msb_decoder  msb_decoder_0
timestamp 1748318706
transform 1 0 0 0 1 400
box 0 0 15596 5868
<< labels >>
flabel metal3 0 0 15596 200 0 FreeSans 256 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 0 400 15596 600 0 FreeSans 256 0 0 0 VDD
port 2 nsew power bidirectional
flabel metal3 5856 13617 10134 13755 0 FreeSans 256 0 0 0 VOUT
port 3 nsew signal bidirectional
flabel metal3 16882 20953 16942 21253 0 FreeSans 256 0 0 0 IN[0]
port 4 nsew signal input
flabel metal3 16756 20953 16816 21253 0 FreeSans 256 0 0 0 IN[1]
port 5 nsew signal input
flabel metal3 16630 20953 16690 21253 0 FreeSans 256 0 0 0 IN[2]
port 6 nsew signal input
flabel metal3 16504 20953 16564 21253 0 FreeSans 256 0 0 0 IN[3]
port 7 nsew signal input
flabel metal3 16378 20953 16438 21253 0 FreeSans 256 0 0 0 IN[4]
port 8 nsew signal input
flabel metal3 16252 20953 16312 21253 0 FreeSans 256 0 0 0 IN[5]
port 9 nsew signal input
flabel metal3 16126 20953 16186 21253 0 FreeSans 256 0 0 0 IN[6]
port 10 nsew signal input
flabel metal3 16000 20953 16060 21253 0 FreeSans 256 0 0 0 IN[7]
port 11 nsew signal input
<< end >>
