magic
tech sky130A
magscale 1 2
timestamp 1748334057
<< dnwell >>
rect 5459 12246 22267 32913
<< nwell >>
rect 5349 32707 22377 33023
rect 5349 12452 5665 32707
rect 22061 12452 22377 32707
rect 5349 12136 22377 12452
<< mvnsubdiff >>
rect 5416 32936 22310 32956
rect 5416 32902 5496 32936
rect 22230 32902 22310 32936
rect 5416 32882 22310 32902
rect 5416 32876 5490 32882
rect 5416 12283 5436 32876
rect 5470 12283 5490 32876
rect 5416 12277 5490 12283
rect 22236 32876 22310 32882
rect 22236 12283 22256 32876
rect 22290 12283 22310 32876
rect 22236 12277 22310 12283
rect 5416 12257 22310 12277
rect 5416 12223 5496 12257
rect 22230 12223 22310 12257
rect 5416 12203 22310 12223
<< mvnsubdiffcont >>
rect 5496 32902 22230 32936
rect 5436 12283 5470 32876
rect 22256 12283 22290 32876
rect 5496 12223 22230 12257
<< locali >>
rect 5436 32902 5496 32936
rect 22230 32902 22290 32936
rect 5436 32876 5470 32902
rect 5436 12257 5470 12283
rect 22256 32876 22290 32902
rect 22256 12257 22290 12283
rect 5436 12223 5496 12257
rect 22230 12223 22290 12257
use toplevel  toplevel_0
timestamp 1748334013
transform 1 0 0 0 1 0
box 0 0 29072 45152
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
