magic
tech sky130A
magscale 1 2
timestamp 1748337984
<< locali >>
rect 150 7240 250 7252
rect 150 6648 156 7240
rect 244 6648 250 7240
rect 150 6636 250 6648
rect 5572 7240 5672 7252
rect 5572 6648 5578 7240
rect 5666 6648 5672 7240
rect 5572 6636 5672 6648
rect 150 6256 253 6268
rect 150 5415 156 6256
rect 244 5415 253 6256
rect 150 5403 253 5415
rect 5572 6256 5672 6268
rect 5572 5415 5578 6256
rect 5666 5415 5672 6256
rect 5572 5403 5672 5415
rect 0 5023 112 5035
rect 0 2373 6 5023
rect 106 2373 112 5023
rect 0 2361 112 2373
rect 5710 5023 5822 5035
rect 5710 2373 5716 5023
rect 5816 2373 5822 5023
rect 5710 2361 5822 2373
rect 150 1981 253 1993
rect 150 1140 156 1981
rect 244 1140 253 1981
rect 150 1128 253 1140
rect 5572 1981 5672 1993
rect 5572 1140 5578 1981
rect 5666 1140 5672 1981
rect 5572 1128 5672 1140
rect 150 748 250 760
rect 150 156 156 748
rect 244 156 250 748
rect 150 144 250 156
rect 5572 748 5672 760
rect 5572 156 5578 748
rect 5666 156 5672 748
rect 5572 144 5672 156
<< viali >>
rect 156 6648 244 7240
rect 5578 6648 5666 7240
rect 156 5415 244 6256
rect 5578 5415 5666 6256
rect 6 2373 106 5023
rect 5716 2373 5816 5023
rect 156 1140 244 1981
rect 5578 1140 5666 1981
rect 156 156 244 748
rect 5578 156 5666 748
<< metal1 >>
rect 0 7240 250 7252
rect 0 6648 6 7240
rect 94 6648 156 7240
rect 244 6648 250 7240
rect 0 6636 250 6648
rect 5572 7240 5822 7252
rect 5572 6648 5578 7240
rect 5666 6648 5728 7240
rect 5816 6648 5822 7240
rect 5572 6636 5822 6648
rect 150 6256 250 6268
rect 150 5415 156 6256
rect 244 5415 250 6256
rect 150 5403 250 5415
rect 5572 6256 5672 6268
rect 5572 5415 5578 6256
rect 5666 5415 5672 6256
rect 5572 5403 5672 5415
rect 0 5023 112 5035
rect 0 2373 6 5023
rect 106 4989 112 5023
rect 5710 5023 5822 5035
rect 5710 4989 5716 5023
rect 106 4808 456 4989
rect 106 4738 386 4808
rect 106 4557 456 4738
rect 552 4808 788 4989
rect 552 4738 635 4808
rect 705 4738 788 4808
rect 552 4557 788 4738
rect 884 4808 1120 4989
rect 884 4738 967 4808
rect 1037 4738 1120 4808
rect 884 4557 1120 4738
rect 1216 4808 1452 4989
rect 1216 4738 1299 4808
rect 1369 4738 1452 4808
rect 1216 4557 1452 4738
rect 1548 4808 1784 4989
rect 1548 4738 1631 4808
rect 1701 4738 1784 4808
rect 1548 4557 1784 4738
rect 1880 4808 2116 4989
rect 1880 4738 1963 4808
rect 2033 4738 2116 4808
rect 1880 4557 2116 4738
rect 2212 4808 2448 4989
rect 2212 4738 2295 4808
rect 2365 4738 2448 4808
rect 2212 4557 2448 4738
rect 2544 4808 2780 4989
rect 2544 4738 2627 4808
rect 2697 4738 2780 4808
rect 2544 4557 2780 4738
rect 106 2839 112 4557
rect 2876 3473 2946 4989
rect 3042 4513 3112 4989
rect 3208 4808 3444 4989
rect 3208 4738 3291 4808
rect 3361 4738 3444 4808
rect 3208 4557 3444 4738
rect 3540 4808 3776 4989
rect 3540 4738 3623 4808
rect 3693 4738 3776 4808
rect 3540 4557 3776 4738
rect 3872 4808 4108 4989
rect 3872 4738 3955 4808
rect 4025 4738 4108 4808
rect 3872 4557 4108 4738
rect 4204 4808 4440 4989
rect 4204 4738 4287 4808
rect 4357 4738 4440 4808
rect 4204 4557 4440 4738
rect 4536 4808 4772 4989
rect 4536 4738 4619 4808
rect 4689 4738 4772 4808
rect 4536 4557 4772 4738
rect 4868 4808 5104 4989
rect 4868 4738 4951 4808
rect 5021 4738 5104 4808
rect 4868 4557 5104 4738
rect 5200 4808 5436 4989
rect 5200 4738 5283 4808
rect 5353 4738 5436 4808
rect 5200 4557 5436 4738
rect 5532 4557 5716 4989
rect 3042 4437 3112 4443
rect 2870 3403 2876 3473
rect 2946 3403 2952 3473
rect 5710 2839 5716 4557
rect 106 2407 290 2839
rect 386 2658 622 2839
rect 386 2588 469 2658
rect 539 2588 622 2658
rect 386 2407 622 2588
rect 718 2658 954 2839
rect 718 2588 801 2658
rect 871 2588 954 2658
rect 718 2407 954 2588
rect 1050 2658 1286 2839
rect 1050 2588 1133 2658
rect 1203 2588 1286 2658
rect 1050 2407 1286 2588
rect 1382 2658 1618 2839
rect 1382 2588 1465 2658
rect 1535 2588 1618 2658
rect 1382 2407 1618 2588
rect 1714 2658 1950 2839
rect 1714 2588 1797 2658
rect 1867 2588 1950 2658
rect 1714 2407 1950 2588
rect 2046 2658 2282 2839
rect 2046 2588 2129 2658
rect 2199 2588 2282 2658
rect 2046 2407 2282 2588
rect 2378 2658 2614 2839
rect 2378 2588 2461 2658
rect 2531 2588 2614 2658
rect 2378 2407 2614 2588
rect 2710 2658 2946 2839
rect 2710 2588 2793 2658
rect 2863 2588 2946 2658
rect 2710 2407 2946 2588
rect 3042 2658 3278 2839
rect 3042 2588 3125 2658
rect 3195 2588 3278 2658
rect 3042 2407 3278 2588
rect 3374 2658 3610 2839
rect 3374 2588 3457 2658
rect 3527 2588 3610 2658
rect 3374 2407 3610 2588
rect 3706 2658 3942 2839
rect 3706 2588 3789 2658
rect 3859 2588 3942 2658
rect 3706 2407 3942 2588
rect 4038 2658 4274 2839
rect 4038 2588 4121 2658
rect 4191 2588 4274 2658
rect 4038 2407 4274 2588
rect 4370 2658 4606 2839
rect 4370 2588 4453 2658
rect 4523 2588 4606 2658
rect 4370 2407 4606 2588
rect 4702 2658 4938 2839
rect 4702 2588 4785 2658
rect 4855 2588 4938 2658
rect 4702 2407 4938 2588
rect 5034 2658 5270 2839
rect 5034 2588 5117 2658
rect 5187 2588 5270 2658
rect 5034 2407 5270 2588
rect 5366 2658 5436 2839
rect 5366 2407 5436 2588
rect 5532 2407 5716 2839
rect 106 2373 112 2407
rect 0 2361 112 2373
rect 5710 2373 5716 2407
rect 5816 2373 5822 5023
rect 5710 2361 5822 2373
rect 150 1981 250 1993
rect 150 1140 156 1981
rect 244 1140 250 1981
rect 150 1128 250 1140
rect 5572 1981 5672 1993
rect 5572 1140 5578 1981
rect 5666 1140 5672 1981
rect 5572 1128 5672 1140
rect 0 748 250 760
rect 0 156 6 748
rect 94 156 156 748
rect 244 156 250 748
rect 0 144 250 156
rect 5572 748 5822 760
rect 5572 156 5578 748
rect 5666 156 5728 748
rect 5816 156 5822 748
rect 5572 144 5822 156
<< via1 >>
rect 6 6648 94 7240
rect 5728 6648 5816 7240
rect 156 5415 244 6256
rect 5578 5415 5666 6256
rect 6 2373 94 5023
rect 386 4738 456 4808
rect 635 4738 705 4808
rect 967 4738 1037 4808
rect 1299 4738 1369 4808
rect 1631 4738 1701 4808
rect 1963 4738 2033 4808
rect 2295 4738 2365 4808
rect 2627 4738 2697 4808
rect 3291 4738 3361 4808
rect 3623 4738 3693 4808
rect 3955 4738 4025 4808
rect 4287 4738 4357 4808
rect 4619 4738 4689 4808
rect 4951 4738 5021 4808
rect 5283 4738 5353 4808
rect 3042 4443 3112 4513
rect 2876 3403 2946 3473
rect 469 2588 539 2658
rect 801 2588 871 2658
rect 1133 2588 1203 2658
rect 1465 2588 1535 2658
rect 1797 2588 1867 2658
rect 2129 2588 2199 2658
rect 2461 2588 2531 2658
rect 2793 2588 2863 2658
rect 3125 2588 3195 2658
rect 3457 2588 3527 2658
rect 3789 2588 3859 2658
rect 4121 2588 4191 2658
rect 4453 2588 4523 2658
rect 4785 2588 4855 2658
rect 5117 2588 5187 2658
rect 5366 2588 5436 2658
rect 5728 2373 5816 5023
rect 156 1140 244 1981
rect 5578 1140 5666 1981
rect 6 156 94 748
rect 5728 156 5816 748
<< metal2 >>
rect 0 7240 100 7396
rect 0 6648 6 7240
rect 94 6648 100 7240
rect 0 5023 100 6648
rect 0 2373 6 5023
rect 94 2373 100 5023
rect 0 748 100 2373
rect 0 156 6 748
rect 94 156 100 748
rect 0 0 100 156
rect 150 6256 250 7396
rect 685 6711 823 7354
rect 961 6883 1099 7021
rect 1237 6883 1375 7021
rect 1513 6883 1651 7021
rect 1789 6883 1927 7021
rect 2065 6883 2203 7021
rect 2341 6883 2479 7021
rect 2617 6883 2755 7021
rect 2893 6883 3031 7021
rect 3169 6883 3307 7021
rect 3445 6883 3583 7021
rect 3721 6883 3859 7021
rect 3997 6883 4135 7021
rect 4273 6883 4411 7021
rect 4549 6883 4687 7021
rect 4825 6883 4963 7021
rect 5101 6883 5239 7021
rect 961 6839 1099 6849
rect 961 6721 971 6839
rect 1089 6721 1099 6839
rect 961 6711 1099 6721
rect 1237 6839 1375 6849
rect 1237 6721 1247 6839
rect 1365 6721 1375 6839
rect 1237 6711 1375 6721
rect 1513 6839 1651 6849
rect 1513 6721 1523 6839
rect 1641 6721 1651 6839
rect 1513 6711 1651 6721
rect 1789 6839 1927 6849
rect 1789 6721 1799 6839
rect 1917 6721 1927 6839
rect 1789 6711 1927 6721
rect 2065 6839 2203 6849
rect 2065 6721 2075 6839
rect 2193 6721 2203 6839
rect 2065 6711 2203 6721
rect 2341 6839 2479 6849
rect 2341 6721 2351 6839
rect 2469 6721 2479 6839
rect 2341 6711 2479 6721
rect 2617 6839 2755 6849
rect 2617 6721 2627 6839
rect 2745 6721 2755 6839
rect 2617 6711 2755 6721
rect 2893 6839 3031 6849
rect 2893 6721 2903 6839
rect 3021 6721 3031 6839
rect 2893 6711 3031 6721
rect 3169 6839 3307 6849
rect 3169 6721 3179 6839
rect 3297 6721 3307 6839
rect 3169 6711 3307 6721
rect 3445 6839 3583 6849
rect 3445 6721 3455 6839
rect 3573 6721 3583 6839
rect 3445 6711 3583 6721
rect 3721 6839 3859 6849
rect 3721 6721 3731 6839
rect 3849 6721 3859 6839
rect 3721 6711 3859 6721
rect 3997 6839 4135 6849
rect 3997 6721 4007 6839
rect 4125 6721 4135 6839
rect 3997 6711 4135 6721
rect 4273 6839 4411 6849
rect 4273 6721 4283 6839
rect 4401 6721 4411 6839
rect 4273 6711 4411 6721
rect 4549 6839 4687 6849
rect 4549 6721 4559 6839
rect 4677 6721 4687 6839
rect 4549 6711 4687 6721
rect 4825 6839 4963 6849
rect 4825 6721 4835 6839
rect 4953 6721 4963 6839
rect 4825 6711 4963 6721
rect 5101 6839 5239 6849
rect 5101 6721 5111 6839
rect 5229 6721 5239 6839
rect 5101 6711 5239 6721
rect 150 5415 156 6256
rect 244 5415 250 6256
rect 5572 6256 5672 7396
rect 583 5704 721 6203
rect 893 6169 963 6178
rect 893 6090 963 6099
rect 1169 6169 1239 6178
rect 1169 6090 1239 6099
rect 1445 6169 1515 6178
rect 1445 6090 1515 6099
rect 1721 6169 1791 6178
rect 1721 6090 1791 6099
rect 1997 6169 2067 6178
rect 1997 6090 2067 6099
rect 2273 6169 2343 6178
rect 2273 6090 2343 6099
rect 2549 6169 2619 6178
rect 2549 6090 2619 6099
rect 2825 6169 2895 6178
rect 2825 6090 2895 6099
rect 3101 6169 3171 6178
rect 3101 6090 3171 6099
rect 3377 6169 3447 6178
rect 3377 6090 3447 6099
rect 3653 6169 3723 6178
rect 3653 6090 3723 6099
rect 3929 6169 3999 6178
rect 3929 6090 3999 6099
rect 4205 6169 4275 6178
rect 4205 6090 4275 6099
rect 4481 6169 4551 6178
rect 4481 6090 4551 6099
rect 4757 6169 4827 6178
rect 4757 6090 4827 6099
rect 5033 6169 5103 6178
rect 5033 6090 5103 6099
rect 150 3468 250 5415
rect 5572 5415 5578 6256
rect 5666 5415 5672 6256
rect 4453 5239 4523 5244
rect 4619 5239 4689 5244
rect 4785 5239 4855 5244
rect 4951 5239 5021 5244
rect 5117 5239 5187 5244
rect 5283 5239 5353 5244
rect 4449 5179 4458 5239
rect 4518 5179 4527 5239
rect 4615 5179 4624 5239
rect 4684 5179 4693 5239
rect 4781 5179 4790 5239
rect 4850 5179 4859 5239
rect 4947 5179 4956 5239
rect 5016 5179 5025 5239
rect 5113 5179 5122 5239
rect 5182 5179 5191 5239
rect 5279 5179 5288 5239
rect 5348 5179 5357 5239
rect 4287 5158 4357 5163
rect 4283 5098 4292 5158
rect 4352 5098 4361 5158
rect 4121 5028 4191 5033
rect 4117 4968 4126 5028
rect 4186 4968 4195 5028
rect 3955 4898 4025 4903
rect 3951 4838 3960 4898
rect 4020 4838 4029 4898
rect 3955 4808 4025 4838
rect 150 3408 155 3468
rect 215 3408 250 3468
rect 150 1981 250 3408
rect 303 4738 386 4808
rect 456 4738 462 4808
rect 629 4738 635 4808
rect 705 4738 711 4808
rect 961 4738 967 4808
rect 1037 4738 1043 4808
rect 1293 4738 1299 4808
rect 1369 4738 1375 4808
rect 1625 4738 1631 4808
rect 1701 4738 1707 4808
rect 1957 4738 1963 4808
rect 2033 4738 2039 4808
rect 2289 4738 2295 4808
rect 2365 4738 2371 4808
rect 2621 4738 2627 4808
rect 2697 4738 2703 4808
rect 3285 4738 3291 4808
rect 3361 4738 3367 4808
rect 3617 4738 3623 4808
rect 3693 4738 3699 4808
rect 3789 4768 3859 4773
rect 303 2217 373 4738
rect 463 2588 469 2658
rect 539 2588 545 2658
rect 469 2217 539 2588
rect 635 2217 705 4738
rect 795 2588 801 2658
rect 871 2588 877 2658
rect 801 2217 871 2588
rect 967 2217 1037 4738
rect 1127 2588 1133 2658
rect 1203 2588 1209 2658
rect 1133 2217 1203 2588
rect 1299 2217 1369 4738
rect 1459 2588 1465 2658
rect 1535 2588 1541 2658
rect 1465 2298 1535 2588
rect 1631 2428 1701 4738
rect 1963 2688 2033 4738
rect 2295 2948 2365 4738
rect 2627 3208 2697 4738
rect 2959 4443 3042 4513
rect 3112 4443 3118 4513
rect 2959 4118 3029 4443
rect 3291 4378 3361 4738
rect 3623 4638 3693 4738
rect 3785 4708 3794 4768
rect 3854 4708 3863 4768
rect 3949 4738 3955 4808
rect 4025 4738 4031 4808
rect 3619 4578 3628 4638
rect 3688 4578 3697 4638
rect 3623 4573 3693 4578
rect 3457 4508 3527 4513
rect 3453 4448 3462 4508
rect 3522 4448 3531 4508
rect 3287 4318 3296 4378
rect 3356 4318 3365 4378
rect 3291 4313 3361 4318
rect 3125 4248 3195 4253
rect 3121 4188 3130 4248
rect 3190 4188 3199 4248
rect 2955 4058 2964 4118
rect 3024 4058 3033 4118
rect 2959 3608 3029 4058
rect 2950 3538 2959 3608
rect 3029 3538 3038 3608
rect 2876 3473 2946 3479
rect 2872 3408 2876 3468
rect 2946 3408 2950 3468
rect 2876 3397 2946 3403
rect 2793 3338 2863 3343
rect 2789 3278 2798 3338
rect 2858 3278 2867 3338
rect 2623 3148 2632 3208
rect 2692 3148 2701 3208
rect 2627 3143 2697 3148
rect 2461 3078 2531 3083
rect 2457 3018 2466 3078
rect 2526 3018 2535 3078
rect 2291 2888 2300 2948
rect 2360 2888 2369 2948
rect 2295 2883 2365 2888
rect 2129 2818 2199 2823
rect 2125 2758 2134 2818
rect 2194 2758 2203 2818
rect 1791 2588 1797 2658
rect 1867 2588 1873 2658
rect 1959 2628 1968 2688
rect 2028 2628 2037 2688
rect 2129 2658 2199 2758
rect 2461 2658 2531 3018
rect 2793 2658 2863 3278
rect 3125 2658 3195 4188
rect 3457 2658 3527 4448
rect 3789 2658 3859 4708
rect 4121 2658 4191 4968
rect 4287 4808 4357 5098
rect 4281 4738 4287 4808
rect 4357 4738 4363 4808
rect 4453 2658 4523 5179
rect 4619 4808 4689 5179
rect 4613 4738 4619 4808
rect 4689 4738 4695 4808
rect 4785 2658 4855 5179
rect 4951 4808 5021 5179
rect 4945 4738 4951 4808
rect 5021 4738 5027 4808
rect 5117 2658 5187 5179
rect 5283 4808 5353 5179
rect 5277 4738 5283 4808
rect 5353 4738 5359 4808
rect 5449 2658 5519 2664
rect 1963 2623 2033 2628
rect 2123 2588 2129 2658
rect 2199 2588 2205 2658
rect 2455 2588 2461 2658
rect 2531 2588 2537 2658
rect 2787 2588 2793 2658
rect 2863 2588 2869 2658
rect 3119 2588 3125 2658
rect 3195 2588 3201 2658
rect 3451 2588 3457 2658
rect 3527 2588 3533 2658
rect 3783 2588 3789 2658
rect 3859 2588 3865 2658
rect 4115 2588 4121 2658
rect 4191 2588 4197 2658
rect 4447 2588 4453 2658
rect 4523 2588 4529 2658
rect 4779 2588 4785 2658
rect 4855 2588 4861 2658
rect 5111 2588 5117 2658
rect 5187 2588 5193 2658
rect 5360 2588 5366 2658
rect 5436 2653 5519 2658
rect 5436 2593 5454 2653
rect 5514 2593 5523 2653
rect 5436 2588 5519 2593
rect 1797 2558 1867 2588
rect 5449 2582 5519 2588
rect 1793 2498 1802 2558
rect 1862 2498 1871 2558
rect 1797 2493 1867 2498
rect 1627 2368 1636 2428
rect 1696 2368 1705 2428
rect 1631 2363 1701 2368
rect 1461 2238 1470 2298
rect 1530 2238 1539 2298
rect 1465 2233 1535 2238
rect 299 2157 308 2217
rect 368 2157 377 2217
rect 465 2157 474 2217
rect 534 2157 543 2217
rect 631 2157 640 2217
rect 700 2157 709 2217
rect 797 2157 806 2217
rect 866 2157 875 2217
rect 963 2157 972 2217
rect 1032 2157 1041 2217
rect 1129 2157 1138 2217
rect 1198 2157 1207 2217
rect 1295 2157 1304 2217
rect 1364 2157 1373 2217
rect 303 2152 373 2157
rect 469 2152 539 2157
rect 635 2152 705 2157
rect 801 2152 871 2157
rect 967 2152 1037 2157
rect 1133 2152 1203 2157
rect 1299 2152 1369 2157
rect 150 1140 156 1981
rect 244 1140 250 1981
rect 5572 1981 5672 5415
rect 719 1297 789 1306
rect 719 1218 789 1227
rect 995 1297 1065 1306
rect 995 1218 1065 1227
rect 1271 1297 1341 1306
rect 1271 1218 1341 1227
rect 1547 1297 1617 1306
rect 1547 1218 1617 1227
rect 1823 1297 1893 1306
rect 1823 1218 1893 1227
rect 2099 1297 2169 1306
rect 2099 1218 2169 1227
rect 2375 1297 2445 1306
rect 2375 1218 2445 1227
rect 2651 1297 2721 1306
rect 2651 1218 2721 1227
rect 2927 1297 2997 1306
rect 2927 1218 2997 1227
rect 3203 1297 3273 1306
rect 3203 1218 3273 1227
rect 3479 1297 3549 1306
rect 3479 1218 3549 1227
rect 3755 1297 3825 1306
rect 3755 1218 3825 1227
rect 4031 1297 4101 1306
rect 4031 1218 4101 1227
rect 4307 1297 4377 1306
rect 4307 1218 4377 1227
rect 4583 1297 4653 1306
rect 4583 1218 4653 1227
rect 4859 1297 4929 1306
rect 4859 1218 4929 1227
rect 5135 1297 5205 1306
rect 5135 1218 5205 1227
rect 150 0 250 1140
rect 5572 1140 5578 1981
rect 5666 1140 5672 1981
rect 583 675 721 685
rect 583 557 593 675
rect 711 557 721 675
rect 583 547 721 557
rect 859 675 997 685
rect 859 557 869 675
rect 987 557 997 675
rect 859 547 997 557
rect 1135 675 1273 685
rect 1135 557 1145 675
rect 1263 557 1273 675
rect 1135 547 1273 557
rect 1411 675 1549 685
rect 1411 557 1421 675
rect 1539 557 1549 675
rect 1411 547 1549 557
rect 1687 675 1825 685
rect 1687 557 1697 675
rect 1815 557 1825 675
rect 1687 547 1825 557
rect 1963 675 2101 685
rect 1963 557 1973 675
rect 2091 557 2101 675
rect 1963 547 2101 557
rect 2239 675 2377 685
rect 2239 557 2249 675
rect 2367 557 2377 675
rect 2239 547 2377 557
rect 2515 675 2653 685
rect 2515 557 2525 675
rect 2643 557 2653 675
rect 2515 547 2653 557
rect 2791 675 2929 685
rect 2791 557 2801 675
rect 2919 557 2929 675
rect 2791 547 2929 557
rect 3067 675 3205 685
rect 3067 557 3077 675
rect 3195 557 3205 675
rect 3067 547 3205 557
rect 3343 675 3481 685
rect 3343 557 3353 675
rect 3471 557 3481 675
rect 3343 547 3481 557
rect 3619 675 3757 685
rect 3619 557 3629 675
rect 3747 557 3757 675
rect 3619 547 3757 557
rect 3895 675 4033 685
rect 3895 557 3905 675
rect 4023 557 4033 675
rect 3895 547 4033 557
rect 4171 675 4309 685
rect 4171 557 4181 675
rect 4299 557 4309 675
rect 4171 547 4309 557
rect 4447 675 4585 685
rect 4447 557 4457 675
rect 4575 557 4585 675
rect 4447 547 4585 557
rect 4723 675 4861 685
rect 4723 557 4733 675
rect 4851 557 4861 675
rect 4723 547 4861 557
rect 4999 675 5137 685
rect 4999 557 5009 675
rect 5127 557 5137 675
rect 4999 547 5137 557
rect 583 375 721 513
rect 859 375 997 513
rect 1135 375 1273 513
rect 1411 375 1549 513
rect 1687 375 1825 513
rect 1963 375 2101 513
rect 2239 375 2377 513
rect 2515 375 2653 513
rect 2791 375 2929 513
rect 3067 375 3205 513
rect 3343 375 3481 513
rect 3619 375 3757 513
rect 3895 375 4033 513
rect 4171 375 4309 513
rect 4447 375 4585 513
rect 4723 375 4861 513
rect 4999 375 5137 513
rect 5572 0 5672 1140
rect 5722 7240 5822 7396
rect 5722 6648 5728 7240
rect 5816 6648 5822 7240
rect 5722 5023 5822 6648
rect 5722 2373 5728 5023
rect 5816 2373 5822 5023
rect 5722 748 5822 2373
rect 5722 156 5728 748
rect 5816 156 5822 748
rect 5722 0 5822 156
<< via2 >>
rect 971 6721 1089 6839
rect 1247 6721 1365 6839
rect 1523 6721 1641 6839
rect 1799 6721 1917 6839
rect 2075 6721 2193 6839
rect 2351 6721 2469 6839
rect 2627 6721 2745 6839
rect 2903 6721 3021 6839
rect 3179 6721 3297 6839
rect 3455 6721 3573 6839
rect 3731 6721 3849 6839
rect 4007 6721 4125 6839
rect 4283 6721 4401 6839
rect 4559 6721 4677 6839
rect 4835 6721 4953 6839
rect 5111 6721 5229 6839
rect 893 6099 963 6169
rect 1169 6099 1239 6169
rect 1445 6099 1515 6169
rect 1721 6099 1791 6169
rect 1997 6099 2067 6169
rect 2273 6099 2343 6169
rect 2549 6099 2619 6169
rect 2825 6099 2895 6169
rect 3101 6099 3171 6169
rect 3377 6099 3447 6169
rect 3653 6099 3723 6169
rect 3929 6099 3999 6169
rect 4205 6099 4275 6169
rect 4481 6099 4551 6169
rect 4757 6099 4827 6169
rect 5033 6099 5103 6169
rect 4458 5179 4518 5239
rect 4624 5179 4684 5239
rect 4790 5179 4850 5239
rect 4956 5179 5016 5239
rect 5122 5179 5182 5239
rect 5288 5179 5348 5239
rect 4292 5098 4352 5158
rect 4126 4968 4186 5028
rect 3960 4838 4020 4898
rect 155 3408 215 3468
rect 3794 4708 3854 4768
rect 3628 4578 3688 4638
rect 3462 4448 3522 4508
rect 3296 4318 3356 4378
rect 3130 4188 3190 4248
rect 2964 4058 3024 4118
rect 2959 3538 3029 3608
rect 2881 3408 2941 3468
rect 2798 3278 2858 3338
rect 2632 3148 2692 3208
rect 2466 3018 2526 3078
rect 2300 2888 2360 2948
rect 2134 2758 2194 2818
rect 1968 2628 2028 2688
rect 5454 2593 5514 2653
rect 1802 2498 1862 2558
rect 1636 2368 1696 2428
rect 1470 2238 1530 2298
rect 308 2157 368 2217
rect 474 2157 534 2217
rect 640 2157 700 2217
rect 806 2157 866 2217
rect 972 2157 1032 2217
rect 1138 2157 1198 2217
rect 1304 2157 1364 2217
rect 719 1227 789 1297
rect 995 1227 1065 1297
rect 1271 1227 1341 1297
rect 1547 1227 1617 1297
rect 1823 1227 1893 1297
rect 2099 1227 2169 1297
rect 2375 1227 2445 1297
rect 2651 1227 2721 1297
rect 2927 1227 2997 1297
rect 3203 1227 3273 1297
rect 3479 1227 3549 1297
rect 3755 1227 3825 1297
rect 4031 1227 4101 1297
rect 4307 1227 4377 1297
rect 4583 1227 4653 1297
rect 4859 1227 4929 1297
rect 5135 1227 5205 1297
rect 593 557 711 675
rect 869 557 987 675
rect 1145 557 1263 675
rect 1421 557 1539 675
rect 1697 557 1815 675
rect 1973 557 2091 675
rect 2249 557 2367 675
rect 2525 557 2643 675
rect 2801 557 2919 675
rect 3077 557 3195 675
rect 3353 557 3471 675
rect 3629 557 3747 675
rect 3905 557 4023 675
rect 4181 557 4299 675
rect 4457 557 4575 675
rect 4733 557 4851 675
rect 5009 557 5127 675
<< metal3 >>
rect 961 6839 5239 6849
rect 961 6721 971 6839
rect 1089 6721 1247 6839
rect 1365 6721 1523 6839
rect 1641 6721 1799 6839
rect 1917 6721 2075 6839
rect 2193 6721 2351 6839
rect 2469 6721 2627 6839
rect 2745 6721 2903 6839
rect 3021 6721 3179 6839
rect 3297 6721 3455 6839
rect 3573 6721 3731 6839
rect 3849 6721 4007 6839
rect 4125 6721 4283 6839
rect 4401 6721 4559 6839
rect 4677 6721 4835 6839
rect 4953 6721 5111 6839
rect 5229 6721 5239 6839
rect 961 6711 5239 6721
rect 5038 6174 5108 6180
rect 888 6169 968 6174
rect 888 6099 893 6169
rect 963 6099 968 6169
rect 888 6094 968 6099
rect 1164 6169 1244 6174
rect 1164 6099 1169 6169
rect 1239 6099 1244 6169
rect 1164 6094 1244 6099
rect 1440 6169 1520 6174
rect 1440 6099 1445 6169
rect 1515 6099 1520 6169
rect 1440 6094 1520 6099
rect 1716 6169 1796 6174
rect 1716 6099 1721 6169
rect 1791 6099 1796 6169
rect 1716 6094 1796 6099
rect 1992 6169 2072 6174
rect 1992 6099 1997 6169
rect 2067 6099 2072 6169
rect 1992 6094 2072 6099
rect 2268 6169 2348 6174
rect 2268 6099 2273 6169
rect 2343 6099 2348 6169
rect 2268 6094 2348 6099
rect 2544 6169 2624 6174
rect 2544 6099 2549 6169
rect 2619 6099 2624 6169
rect 2544 6094 2624 6099
rect 2820 6169 2900 6174
rect 2820 6099 2825 6169
rect 2895 6099 2900 6169
rect 2820 6094 2900 6099
rect 3096 6169 3176 6174
rect 3096 6099 3101 6169
rect 3171 6099 3176 6169
rect 3096 6094 3176 6099
rect 3372 6169 3452 6174
rect 3372 6099 3377 6169
rect 3447 6099 3452 6169
rect 3372 6094 3452 6099
rect 3648 6169 3728 6174
rect 3648 6099 3653 6169
rect 3723 6099 3728 6169
rect 3648 6094 3728 6099
rect 3924 6169 4004 6174
rect 3924 6099 3929 6169
rect 3999 6099 4004 6169
rect 3924 6094 4004 6099
rect 4200 6169 4280 6174
rect 4200 6099 4205 6169
rect 4275 6099 4280 6169
rect 4200 6094 4280 6099
rect 4476 6169 4556 6174
rect 4476 6099 4481 6169
rect 4551 6099 4556 6169
rect 4476 6094 4556 6099
rect 4752 6169 4832 6174
rect 4752 6099 4757 6169
rect 4827 6099 4832 6169
rect 4752 6094 4832 6099
rect 5028 6169 5108 6174
rect 5028 6099 5033 6169
rect 5103 6099 5108 6169
rect 5028 6094 5108 6099
rect 893 4123 963 6094
rect 1169 4253 1239 6094
rect 1445 4383 1515 6094
rect 1721 4513 1791 6094
rect 1997 4643 2067 6094
rect 2273 4773 2343 6094
rect 2549 4903 2619 6094
rect 2825 5033 2895 6094
rect 3101 5163 3171 6094
rect 3377 5293 3447 6094
rect 3653 5423 3723 6094
rect 3929 5553 3999 6094
rect 4205 5683 4275 6094
rect 4481 5813 4551 6094
rect 4757 5943 4827 6094
rect 5033 6078 5108 6094
rect 5033 6008 5519 6078
rect 4757 5873 5353 5943
rect 4481 5743 5187 5813
rect 4205 5613 5021 5683
rect 3929 5483 4855 5553
rect 3653 5353 4689 5423
rect 3377 5239 4523 5293
rect 3377 5223 4458 5239
rect 4453 5179 4458 5223
rect 4518 5179 4523 5239
rect 4453 5174 4523 5179
rect 4619 5239 4689 5353
rect 4619 5179 4624 5239
rect 4684 5179 4689 5239
rect 4619 5174 4689 5179
rect 4785 5239 4855 5483
rect 4785 5179 4790 5239
rect 4850 5179 4855 5239
rect 4785 5174 4855 5179
rect 4951 5239 5021 5613
rect 4951 5179 4956 5239
rect 5016 5179 5021 5239
rect 4951 5174 5021 5179
rect 5117 5239 5187 5743
rect 5117 5179 5122 5239
rect 5182 5179 5187 5239
rect 5117 5174 5187 5179
rect 5283 5239 5353 5873
rect 5283 5179 5288 5239
rect 5348 5179 5353 5239
rect 5283 5174 5353 5179
rect 3101 5158 4357 5163
rect 3101 5098 4292 5158
rect 4352 5098 4357 5158
rect 3101 5093 4357 5098
rect 2825 5028 4191 5033
rect 2825 4968 4126 5028
rect 4186 4968 4191 5028
rect 2825 4963 4191 4968
rect 2549 4898 4025 4903
rect 2549 4838 3960 4898
rect 4020 4838 4025 4898
rect 2549 4833 4025 4838
rect 2273 4768 3859 4773
rect 2273 4708 3794 4768
rect 3854 4708 3859 4768
rect 2273 4703 3859 4708
rect 1997 4638 3693 4643
rect 1997 4578 3628 4638
rect 3688 4578 3693 4638
rect 1997 4573 3693 4578
rect 1721 4508 3527 4513
rect 1721 4448 3462 4508
rect 3522 4448 3527 4508
rect 1721 4443 3527 4448
rect 1445 4378 3361 4383
rect 1445 4318 3296 4378
rect 3356 4318 3361 4378
rect 1445 4313 3361 4318
rect 1169 4248 3195 4253
rect 1169 4188 3130 4248
rect 3190 4188 3195 4248
rect 1169 4183 3195 4188
rect 893 4118 3029 4123
rect 893 4058 2964 4118
rect 3024 4058 3029 4118
rect 893 4053 3029 4058
rect 2954 3608 3034 3613
rect 2954 3538 2959 3608
rect 3029 3538 5340 3608
rect 2954 3533 3034 3538
rect 150 3468 5205 3473
rect 150 3408 155 3468
rect 215 3408 2881 3468
rect 2941 3408 5205 3468
rect 150 3403 5205 3408
rect 2793 3338 4929 3343
rect 2793 3278 2798 3338
rect 2858 3278 4929 3338
rect 2793 3273 4929 3278
rect 2627 3208 4653 3213
rect 2627 3148 2632 3208
rect 2692 3148 4653 3208
rect 2627 3143 4653 3148
rect 2461 3078 4377 3083
rect 2461 3018 2466 3078
rect 2526 3018 4377 3078
rect 2461 3013 4377 3018
rect 2295 2948 4101 2953
rect 2295 2888 2300 2948
rect 2360 2888 4101 2948
rect 2295 2883 4101 2888
rect 2129 2818 3825 2823
rect 2129 2758 2134 2818
rect 2194 2758 3825 2818
rect 2129 2753 3825 2758
rect 1963 2688 3549 2693
rect 1963 2628 1968 2688
rect 2028 2628 3549 2688
rect 1963 2623 3549 2628
rect 1797 2558 3273 2563
rect 1797 2498 1802 2558
rect 1862 2498 3273 2558
rect 1797 2493 3273 2498
rect 1631 2428 2997 2433
rect 1631 2368 1636 2428
rect 1696 2368 2997 2428
rect 1631 2363 2997 2368
rect 1465 2298 2721 2303
rect 1465 2238 1470 2298
rect 1530 2238 2721 2298
rect 1465 2233 2721 2238
rect 303 2217 373 2222
rect 303 2157 308 2217
rect 368 2157 373 2217
rect 303 1388 373 2157
rect 469 2217 539 2222
rect 469 2157 474 2217
rect 534 2157 539 2217
rect 469 1523 539 2157
rect 635 2217 705 2222
rect 635 2157 640 2217
rect 700 2157 705 2217
rect 635 1653 705 2157
rect 801 2217 871 2222
rect 801 2157 806 2217
rect 866 2157 871 2217
rect 801 1783 871 2157
rect 967 2217 1037 2222
rect 967 2157 972 2217
rect 1032 2157 1037 2217
rect 967 1913 1037 2157
rect 1133 2217 1203 2222
rect 1133 2157 1138 2217
rect 1198 2157 1203 2217
rect 1133 2043 1203 2157
rect 1299 2217 1369 2222
rect 1299 2157 1304 2217
rect 1364 2173 1369 2217
rect 1364 2157 2445 2173
rect 1299 2103 2445 2157
rect 1133 1973 2169 2043
rect 967 1843 1893 1913
rect 801 1713 1617 1783
rect 635 1583 1341 1653
rect 469 1453 1065 1523
rect 303 1318 789 1388
rect 714 1302 789 1318
rect 995 1302 1065 1453
rect 1271 1302 1341 1583
rect 1547 1302 1617 1713
rect 1823 1302 1893 1843
rect 2099 1302 2169 1973
rect 2375 1302 2445 2103
rect 2651 1302 2721 2233
rect 2927 1302 2997 2363
rect 3203 1302 3273 2493
rect 3479 1302 3549 2623
rect 3755 1302 3825 2753
rect 4031 1302 4101 2883
rect 4307 1302 4377 3013
rect 4583 1302 4653 3143
rect 4859 1302 4929 3273
rect 5135 1302 5205 3403
rect 714 1297 794 1302
rect 714 1227 719 1297
rect 789 1227 794 1297
rect 714 1222 794 1227
rect 990 1297 1070 1302
rect 990 1227 995 1297
rect 1065 1227 1070 1297
rect 990 1222 1070 1227
rect 1266 1297 1346 1302
rect 1266 1227 1271 1297
rect 1341 1227 1346 1297
rect 1266 1222 1346 1227
rect 1542 1297 1622 1302
rect 1542 1227 1547 1297
rect 1617 1227 1622 1297
rect 1542 1222 1622 1227
rect 1818 1297 1898 1302
rect 1818 1227 1823 1297
rect 1893 1227 1898 1297
rect 1818 1222 1898 1227
rect 2094 1297 2174 1302
rect 2094 1227 2099 1297
rect 2169 1227 2174 1297
rect 2094 1222 2174 1227
rect 2370 1297 2450 1302
rect 2370 1227 2375 1297
rect 2445 1227 2450 1297
rect 2370 1222 2450 1227
rect 2646 1297 2726 1302
rect 2646 1227 2651 1297
rect 2721 1227 2726 1297
rect 2646 1222 2726 1227
rect 2922 1297 3002 1302
rect 2922 1227 2927 1297
rect 2997 1227 3002 1297
rect 2922 1222 3002 1227
rect 3198 1297 3278 1302
rect 3198 1227 3203 1297
rect 3273 1227 3278 1297
rect 3198 1222 3278 1227
rect 3474 1297 3554 1302
rect 3474 1227 3479 1297
rect 3549 1227 3554 1297
rect 3474 1222 3554 1227
rect 3750 1297 3830 1302
rect 3750 1227 3755 1297
rect 3825 1227 3830 1297
rect 3750 1222 3830 1227
rect 4026 1297 4106 1302
rect 4026 1227 4031 1297
rect 4101 1227 4106 1297
rect 4026 1222 4106 1227
rect 4302 1297 4382 1302
rect 4302 1227 4307 1297
rect 4377 1227 4382 1297
rect 4302 1222 4382 1227
rect 4578 1297 4658 1302
rect 4578 1227 4583 1297
rect 4653 1227 4658 1297
rect 4578 1222 4658 1227
rect 4854 1297 4934 1302
rect 4854 1227 4859 1297
rect 4929 1227 4934 1297
rect 4854 1222 4934 1227
rect 5130 1297 5210 1302
rect 5130 1227 5135 1297
rect 5205 1227 5210 1297
rect 5130 1222 5210 1227
rect 5270 815 5340 3538
rect 5449 2663 5519 6008
rect 5444 2653 5524 2663
rect 5444 2593 5454 2653
rect 5514 2593 5524 2653
rect 5444 2583 5524 2593
rect 893 745 5340 815
rect 893 685 963 745
rect 1445 685 1515 745
rect 1997 685 2067 745
rect 2549 685 2619 745
rect 3101 685 3171 745
rect 3653 685 3723 745
rect 4205 685 4275 745
rect 4757 685 4827 745
rect 583 675 721 685
rect 583 557 593 675
rect 711 557 721 675
rect 583 547 721 557
rect 859 675 997 685
rect 859 557 869 675
rect 987 557 997 675
rect 859 547 997 557
rect 1135 675 1273 685
rect 1135 557 1145 675
rect 1263 557 1273 675
rect 1135 547 1273 557
rect 1411 675 1549 685
rect 1411 557 1421 675
rect 1539 557 1549 675
rect 1411 547 1549 557
rect 1687 675 1825 685
rect 1687 557 1697 675
rect 1815 557 1825 675
rect 1687 547 1825 557
rect 1963 675 2101 685
rect 1963 557 1973 675
rect 2091 557 2101 675
rect 1963 547 2101 557
rect 2239 675 2377 685
rect 2239 557 2249 675
rect 2367 557 2377 675
rect 2239 547 2377 557
rect 2515 675 2653 685
rect 2515 557 2525 675
rect 2643 557 2653 675
rect 2515 547 2653 557
rect 2791 675 2929 685
rect 2791 557 2801 675
rect 2919 557 2929 675
rect 2791 547 2929 557
rect 3067 675 3205 685
rect 3067 557 3077 675
rect 3195 557 3205 675
rect 3067 547 3205 557
rect 3343 675 3481 685
rect 3343 557 3353 675
rect 3471 557 3481 675
rect 3343 547 3481 557
rect 3619 675 3757 685
rect 3619 557 3629 675
rect 3747 557 3757 675
rect 3619 547 3757 557
rect 3895 675 4033 685
rect 3895 557 3905 675
rect 4023 557 4033 675
rect 3895 547 4033 557
rect 4171 675 4309 685
rect 4171 557 4181 675
rect 4299 557 4309 675
rect 4171 547 4309 557
rect 4447 675 4585 685
rect 4447 557 4457 675
rect 4575 557 4585 675
rect 4447 547 4585 557
rect 4723 675 4861 685
rect 4723 557 4733 675
rect 4851 557 4861 675
rect 4723 547 4861 557
rect 4999 675 5137 685
rect 4999 557 5009 675
rect 5127 557 5137 675
rect 4999 547 5137 557
rect 617 487 687 547
rect 1169 487 1239 547
rect 1721 487 1791 547
rect 2273 487 2343 547
rect 2825 487 2895 547
rect 3377 487 3447 547
rect 3929 487 3999 547
rect 4481 487 4551 547
rect 5033 487 5103 547
rect 5449 487 5519 2583
rect 617 417 5519 487
use passgates  passgates_0
timestamp 1748309517
transform -1 0 5681 0 -1 7396
box 0 0 5540 2076
use passgates  passgates_2
timestamp 1748309517
transform 1 0 141 0 1 0
box 0 0 5540 2076
use sky130_fd_pr__res_xhigh_po_0p35_7C4M5Y  sky130_fd_pr__res_xhigh_po_0p35_7C4M5Y_0
timestamp 1748333645
transform 1 0 2911 0 1 3698
box -2911 -1511 2911 1511
<< labels >>
flabel metal2 0 0 100 7214 1 FreeSans 400 0 0 0 VSS
port 1 n ground bidirectional
flabel metal2 150 0 250 7214 1 FreeSans 400 0 0 0 VDD
port 2 n power bidirectional
flabel metal3 617 417 5519 487 1 FreeSans 400 0 0 0 A
flabel metal3 893 745 5340 815 1 FreeSans 400 0 0 0 B
flabel metal2 583 375 721 513 1 FreeSans 400 0 0 0 C[0]
port 20 n signal default
flabel metal2 859 375 997 513 1 FreeSans 400 0 0 0 C[1]
port 21 n signal default
flabel metal2 1135 375 1273 513 1 FreeSans 400 0 0 0 C[2]
port 22 n signal default
flabel metal2 1411 375 1549 513 1 FreeSans 400 0 0 0 C[3]
port 23 n signal default
flabel metal2 1687 375 1825 513 1 FreeSans 400 0 0 0 C[4]
port 24 n signal default
flabel metal2 1963 375 2101 513 1 FreeSans 400 0 0 0 C[5]
port 25 n signal default
flabel metal2 2239 375 2377 513 1 FreeSans 400 0 0 0 C[6]
port 26 n signal default
flabel metal2 2515 375 2653 513 1 FreeSans 400 0 0 0 C[7]
port 27 n signal default
flabel metal2 2791 375 2929 513 1 FreeSans 400 0 0 0 C[8]
port 28 n signal default
flabel metal2 3067 375 3205 513 1 FreeSans 400 0 0 0 C[9]
port 29 n signal default
flabel metal2 3343 375 3481 513 1 FreeSans 400 0 0 0 C[10]
port 30 n signal default
flabel metal2 3619 375 3757 513 1 FreeSans 400 0 0 0 C[11]
port 31 n signal default
flabel metal2 3895 375 4033 513 1 FreeSans 400 0 0 0 C[12]
port 32 n signal default
flabel metal2 4171 375 4309 513 1 FreeSans 400 0 0 0 C[13]
port 33 n signal default
flabel metal2 4447 375 4585 513 1 FreeSans 400 0 0 0 C[14]
port 34 n signal default
flabel metal2 4723 375 4861 513 1 FreeSans 400 0 0 0 C[15]
port 35 n signal default
flabel metal2 4999 375 5137 513 1 FreeSans 400 0 0 0 C[16]
port 36 n signal default
flabel metal3 961 6711 5239 6849 1 FreeSans 400 0 0 0 VOUT
port 3 n signal default
flabel metal2 5101 6883 5239 7021 1 FreeSans 400 0 0 0 D[0]
port 4 n signal default
flabel metal2 4825 6883 4963 7021 1 FreeSans 400 0 0 0 D[1]
port 5 n signal default
flabel metal2 4549 6883 4687 7021 1 FreeSans 400 0 0 0 D[2]
port 6 n signal default
flabel metal2 4273 6883 4411 7021 1 FreeSans 400 0 0 0 D[3]
port 7 n signal default
flabel metal2 3997 6883 4135 7021 1 FreeSans 400 0 0 0 D[4]
port 8 n signal default
flabel metal2 3721 6883 3859 7021 1 FreeSans 400 0 0 0 D[5]
port 9 n signal default
flabel metal2 3445 6883 3583 7021 1 FreeSans 400 0 0 0 D[6]
port 10 n signal default
flabel metal2 3169 6883 3307 7021 1 FreeSans 400 0 0 0 D[7]
port 11 n signal default
flabel metal2 2893 6883 3031 7021 1 FreeSans 400 0 0 0 D[8]
port 12 n signal default
flabel metal2 2617 6883 2755 7021 1 FreeSans 400 0 0 0 D[9]
port 13 n signal default
flabel metal2 2341 6883 2479 7021 1 FreeSans 400 0 0 0 D[10]
port 14 n signal default
flabel metal2 2065 6883 2203 7021 1 FreeSans 400 0 0 0 D[11]
port 15 n signal default
flabel metal2 1789 6883 1927 7021 1 FreeSans 400 0 0 0 D[12]
port 16 n signal default
flabel metal2 1513 6883 1651 7021 1 FreeSans 400 0 0 0 D[13]
port 17 n signal default
flabel metal2 1237 6883 1375 7021 1 FreeSans 400 0 0 0 D[14]
port 18 n signal default
flabel metal2 961 6883 1099 7021 1 FreeSans 400 0 0 0 D[15]
port 19 n signal default
<< end >>
