magic
tech sky130A
magscale 1 2
timestamp 1748060222
<< metal1 >>
rect -166 12648 -160 12700
rect -108 12648 -102 12700
rect -243 11306 -237 11358
rect -185 11306 -179 11358
rect -228 8674 -194 11306
rect -151 10016 -117 12648
rect 65 10945 71 10997
rect 123 10945 129 10997
rect -166 9964 -160 10016
rect -108 9964 -102 10016
rect -243 8622 -237 8674
rect -185 8622 -179 8674
rect -228 5990 -194 8622
rect -151 7338 -117 9964
rect -12 8261 -6 8313
rect 46 8261 52 8313
rect -160 7332 -108 7338
rect -160 7274 -108 7280
rect -243 5938 -237 5990
rect -185 5938 -179 5990
rect -228 3306 -194 5938
rect -151 4648 -117 7274
rect -89 5577 -83 5629
rect -31 5577 -25 5629
rect -166 4596 -160 4648
rect -108 4596 -102 4648
rect -243 3254 -237 3306
rect -185 3254 -179 3306
rect -166 2893 -160 2945
rect -108 2893 -102 2945
rect -151 1319 -117 2893
rect -166 1267 -160 1319
rect -108 1267 -102 1319
rect -74 706 -40 5577
rect 3 2661 37 8261
rect -12 2609 -6 2661
rect 46 2609 52 2661
rect 80 2048 114 10945
rect 65 1996 71 2048
rect 123 1996 129 2048
rect -89 654 -83 706
rect -31 654 -25 706
<< via1 >>
rect -160 12648 -108 12700
rect -237 11306 -185 11358
rect 71 10945 123 10997
rect -160 9964 -108 10016
rect -237 8622 -185 8674
rect -6 8261 46 8313
rect -160 7280 -108 7332
rect -237 5938 -185 5990
rect -83 5577 -31 5629
rect -160 4596 -108 4648
rect -237 3254 -185 3306
rect -160 2893 -108 2945
rect -160 1267 -108 1319
rect -6 2609 46 2661
rect 71 1996 123 2048
rect -83 654 -31 706
<< metal2 >>
rect 1859 13401 1919 13410
rect 1919 13354 2918 13388
rect 1859 13332 1919 13341
rect -160 12700 -108 12706
rect -108 12657 315 12691
rect 2772 12657 2918 12691
rect -160 12642 -108 12648
rect 1859 12059 1919 12068
rect 1919 12012 2918 12046
rect 1859 11990 1919 11999
rect -237 11358 -185 11364
rect -185 11315 315 11349
rect 2772 11315 2918 11349
rect -237 11300 -185 11306
rect 71 10997 123 11003
rect 123 10954 272 10988
rect 71 10939 123 10945
rect 1859 10717 1919 10726
rect 1919 10670 2918 10704
rect 1859 10648 1919 10657
rect -160 10016 -108 10022
rect -108 9973 315 10007
rect 2772 9973 2918 10007
rect -160 9958 -108 9964
rect 1859 9375 1919 9384
rect 1919 9328 2918 9362
rect 1859 9306 1919 9315
rect -237 8674 -185 8680
rect -185 8631 315 8665
rect 2772 8631 2918 8665
rect -237 8616 -185 8622
rect -6 8313 46 8319
rect 46 8270 272 8304
rect -6 8255 46 8261
rect 1859 8033 1919 8042
rect 1919 7986 2918 8020
rect 1859 7964 1919 7973
rect -166 7280 -160 7332
rect -108 7323 -102 7332
rect -108 7289 315 7323
rect 2772 7289 2918 7323
rect -108 7280 -102 7289
rect 1859 6691 1919 6700
rect 1919 6644 2918 6678
rect 1859 6622 1919 6631
rect -237 5990 -185 5996
rect -185 5947 315 5981
rect 2772 5947 2918 5981
rect -237 5932 -185 5938
rect -83 5629 -31 5635
rect -31 5586 272 5620
rect -83 5571 -31 5577
rect 1859 5349 1919 5358
rect 1919 5302 2918 5336
rect 1859 5280 1919 5289
rect -160 4648 -108 4654
rect -305 4605 -160 4639
rect -108 4605 572 4639
rect 2772 4605 2918 4639
rect -160 4590 -108 4596
rect 1859 4007 1919 4016
rect 1919 3960 2918 3994
rect 1859 3938 1919 3947
rect -237 3306 -185 3312
rect -305 3263 -237 3297
rect -185 3263 572 3297
rect 2772 3263 2918 3297
rect -237 3248 -185 3254
rect -160 2945 -108 2951
rect -108 2902 272 2936
rect -160 2887 -108 2893
rect -6 2661 46 2667
rect 1859 2665 1919 2674
rect 46 2618 1859 2652
rect -6 2603 46 2609
rect 1859 2596 1919 2605
rect 71 2048 123 2054
rect 123 2005 2206 2039
rect 71 1990 123 1996
rect -305 1921 572 1955
rect 2172 1921 2206 2005
rect -160 1319 -108 1325
rect 1859 1323 1919 1332
rect -108 1276 1859 1310
rect -160 1261 -108 1267
rect 1859 1254 1919 1263
rect -83 706 -31 712
rect -31 663 2206 697
rect -83 648 -31 654
rect -305 579 572 613
rect 2172 579 2206 663
rect 148 218 272 252
<< via2 >>
rect 1859 13341 1919 13401
rect 1859 11999 1919 12059
rect 1859 10657 1919 10717
rect 1859 9315 1919 9375
rect 1859 7973 1919 8033
rect 1859 6631 1919 6691
rect 1859 5289 1919 5349
rect 1859 3947 1919 4007
rect 1859 2605 1919 2665
rect 1859 1263 1919 1323
<< metal3 >>
rect 1854 13401 1924 13406
rect 1854 13341 1859 13401
rect 1919 13341 1924 13401
rect 1854 13336 1924 13341
rect 209 36 269 13304
rect 509 36 569 13304
rect 809 36 869 13304
rect 1109 36 1169 13304
rect 1409 36 1469 13304
rect 1709 36 1769 13304
rect 1859 12540 1919 13336
rect 1854 12059 1924 12064
rect 1854 11999 1859 12059
rect 1919 11999 1924 12059
rect 1854 11994 1924 11999
rect 1859 11198 1919 11994
rect 1854 10717 1924 10722
rect 1854 10657 1859 10717
rect 1919 10657 1924 10717
rect 1854 10652 1924 10657
rect 1859 9856 1919 10652
rect 1854 9375 1924 9380
rect 1854 9315 1859 9375
rect 1919 9315 1924 9375
rect 1854 9310 1924 9315
rect 1859 8514 1919 9310
rect 1854 8033 1924 8038
rect 1854 7973 1859 8033
rect 1919 7973 1924 8033
rect 1854 7968 1924 7973
rect 1859 7172 1919 7968
rect 1854 6691 1924 6696
rect 1854 6631 1859 6691
rect 1919 6631 1924 6691
rect 1854 6626 1924 6631
rect 1859 5830 1919 6626
rect 1854 5349 1924 5354
rect 1854 5289 1859 5349
rect 1919 5289 1924 5349
rect 1854 5284 1924 5289
rect 1859 4488 1919 5284
rect 1854 4007 1924 4012
rect 1854 3947 1859 4007
rect 1919 3947 1924 4007
rect 1854 3942 1924 3947
rect 1859 3146 1919 3942
rect 1854 2665 1924 2670
rect 1854 2605 1859 2665
rect 1919 2605 1924 2665
rect 1854 2600 1924 2605
rect 1859 1804 1919 2600
rect 1854 1323 1924 1328
rect 1854 1263 1859 1323
rect 1919 1263 1924 1323
rect 1854 1258 1924 1263
rect 1859 462 1919 1258
rect 2009 36 2069 13304
rect 2309 36 2369 13304
rect 2609 36 2669 13304
use decoder2  x1
array 0 0 2996 0 4 2684
timestamp 1748060222
transform 1 0 0 0 1 0
box 0 0 2996 2634
<< labels >>
flabel metal3 209 36 269 13304 0 FreeSans 128 0 0 0 VDD
port 0 nsew
flabel metal3 509 36 569 13304 0 FreeSans 128 0 0 0 VSS
port 21 nsew
flabel metal2 -305 579 572 613 0 FreeSans 128 0 0 0 D[2]
port 7 nsew
flabel metal2 -305 1921 572 1955 0 FreeSans 128 0 0 0 D[3]
port 13 nsew
flabel metal2 -305 3263 572 3297 0 FreeSans 128 0 0 0 D[0]
port 11 nsew
flabel metal2 -305 4605 572 4639 0 FreeSans 128 0 0 0 D[1]
port 9 nsew
flabel metal2 2772 3960 2918 3994 0 FreeSans 128 0 0 0 U[0]
port 10 nsew
flabel metal2 2772 3263 2918 3297 0 FreeSans 128 0 0 0 U[1]
port 6 nsew
flabel metal2 2772 5302 2918 5336 0 FreeSans 128 0 0 0 U[2]
port 4 nsew
flabel metal2 2772 4605 2918 4639 0 FreeSans 128 0 0 0 U[3]
port 2 nsew
flabel metal2 2772 6644 2918 6678 0 FreeSans 128 0 0 0 U[4]
port 20 nsew
flabel metal2 2772 5947 2918 5981 0 FreeSans 128 0 0 0 U[5]
port 18 nsew
flabel metal2 2772 7986 2918 8020 0 FreeSans 128 0 0 0 U[6]
port 16 nsew
flabel metal2 2772 7289 2918 7323 0 FreeSans 128 0 0 0 U[7]
port 14 nsew
flabel metal2 2772 9328 2918 9362 0 FreeSans 128 0 0 0 U[8]
port 8 nsew
flabel metal2 2772 8631 2918 8665 0 FreeSans 128 0 0 0 U[9]
port 5 nsew
flabel metal2 2772 10670 2918 10704 0 FreeSans 128 0 0 0 U[10]
port 3 nsew
flabel metal2 2772 9973 2918 10007 0 FreeSans 128 0 0 0 U[11]
port 1 nsew
flabel metal2 2772 12012 2918 12046 0 FreeSans 128 0 0 0 U[12]
port 19 nsew
flabel metal2 2772 11315 2918 11349 0 FreeSans 128 0 0 0 U[13]
port 17 nsew
flabel metal2 2772 13354 2918 13388 0 FreeSans 128 0 0 0 U[14]
port 15 nsew
flabel metal2 2772 12657 2918 12691 0 FreeSans 128 0 0 0 U[15]
port 12 nsew
flabel metal2 148 218 272 252 1 FreeSans 400 0 0 0 EN
port 22 n signal input
<< end >>
